

module mnist_model
(
  input CLK,
  input RESETN,
  output reg irq,
  output reg [32-1:0] maxi_awaddr,
  output reg [8-1:0] maxi_awlen,
  output [3-1:0] maxi_awsize,
  output [2-1:0] maxi_awburst,
  output [1-1:0] maxi_awlock,
  output [4-1:0] maxi_awcache,
  output [3-1:0] maxi_awprot,
  output [4-1:0] maxi_awqos,
  output [2-1:0] maxi_awuser,
  output reg maxi_awvalid,
  input maxi_awready,
  output [32-1:0] maxi_wdata,
  output [4-1:0] maxi_wstrb,
  output maxi_wlast,
  output maxi_wvalid,
  input maxi_wready,
  input [2-1:0] maxi_bresp,
  input maxi_bvalid,
  output maxi_bready,
  output reg [32-1:0] maxi_araddr,
  output reg [8-1:0] maxi_arlen,
  output [3-1:0] maxi_arsize,
  output [2-1:0] maxi_arburst,
  output [1-1:0] maxi_arlock,
  output [4-1:0] maxi_arcache,
  output [3-1:0] maxi_arprot,
  output [4-1:0] maxi_arqos,
  output [2-1:0] maxi_aruser,
  output reg maxi_arvalid,
  input maxi_arready,
  input [32-1:0] maxi_rdata,
  input [2-1:0] maxi_rresp,
  input maxi_rlast,
  input maxi_rvalid,
  output maxi_rready,
  input [32-1:0] saxi_awaddr,
  input [4-1:0] saxi_awcache,
  input [3-1:0] saxi_awprot,
  input saxi_awvalid,
  output saxi_awready,
  input [32-1:0] saxi_wdata,
  input [4-1:0] saxi_wstrb,
  input saxi_wvalid,
  output saxi_wready,
  output [2-1:0] saxi_bresp,
  output reg saxi_bvalid,
  input saxi_bready,
  input [32-1:0] saxi_araddr,
  input [4-1:0] saxi_arcache,
  input [3-1:0] saxi_arprot,
  input saxi_arvalid,
  output saxi_arready,
  output reg [32-1:0] saxi_rdata,
  output [2-1:0] saxi_rresp,
  output reg saxi_rvalid,
  input saxi_rready
);

  wire RESETN_inv;
  assign RESETN_inv = !RESETN;
  wire RESETN_inv_buf;
  reg _RESETN_inv_1;
  reg _RESETN_inv_2;
  assign RESETN_inv_buf = _RESETN_inv_2;
  assign maxi_awsize = 2;
  assign maxi_awburst = 1;
  assign maxi_awlock = 0;
  assign maxi_awcache = 3;
  assign maxi_awprot = 0;
  assign maxi_awqos = 0;
  assign maxi_awuser = 0;
  reg [32-1:0] _maxi_wdata_sb_0;
  reg [4-1:0] _maxi_wstrb_sb_0;
  reg _maxi_wlast_sb_0;
  reg _maxi_wvalid_sb_0;
  wire _maxi_wready_sb_0;
  wire _sb_maxi_writedata_s_value_0;
  assign _sb_maxi_writedata_s_value_0 = _maxi_wlast_sb_0;
  wire [4-1:0] _sb_maxi_writedata_s_value_1;
  assign _sb_maxi_writedata_s_value_1 = _maxi_wstrb_sb_0;
  wire [32-1:0] _sb_maxi_writedata_s_value_2;
  assign _sb_maxi_writedata_s_value_2 = _maxi_wdata_sb_0;
  wire [37-1:0] _sb_maxi_writedata_s_data_3;
  assign _sb_maxi_writedata_s_data_3 = { _sb_maxi_writedata_s_value_0, _sb_maxi_writedata_s_value_1, _sb_maxi_writedata_s_value_2 };
  wire _sb_maxi_writedata_s_valid_4;
  assign _sb_maxi_writedata_s_valid_4 = _maxi_wvalid_sb_0;
  wire _sb_maxi_writedata_m_ready_5;
  assign _sb_maxi_writedata_m_ready_5 = maxi_wready;
  reg [37-1:0] _sb_maxi_writedata_data_6;
  reg _sb_maxi_writedata_valid_7;
  wire _sb_maxi_writedata_ready_8;
  reg [37-1:0] _sb_maxi_writedata_tmp_data_9;
  reg _sb_maxi_writedata_tmp_valid_10;
  wire [37-1:0] _sb_maxi_writedata_next_data_11;
  wire _sb_maxi_writedata_next_valid_12;
  assign _sb_maxi_writedata_ready_8 = !_sb_maxi_writedata_tmp_valid_10;
  assign _sb_maxi_writedata_next_data_11 = (_sb_maxi_writedata_tmp_valid_10)? _sb_maxi_writedata_tmp_data_9 : _sb_maxi_writedata_s_data_3;
  assign _sb_maxi_writedata_next_valid_12 = _sb_maxi_writedata_tmp_valid_10 || _sb_maxi_writedata_s_valid_4;
  wire _sb_maxi_writedata_m_value_13;
  assign _sb_maxi_writedata_m_value_13 = _sb_maxi_writedata_data_6[36:36];
  wire [4-1:0] _sb_maxi_writedata_m_value_14;
  assign _sb_maxi_writedata_m_value_14 = _sb_maxi_writedata_data_6[35:32];
  wire [32-1:0] _sb_maxi_writedata_m_value_15;
  assign _sb_maxi_writedata_m_value_15 = _sb_maxi_writedata_data_6[31:0];
  assign _maxi_wready_sb_0 = _sb_maxi_writedata_ready_8;
  assign maxi_wdata = _sb_maxi_writedata_m_value_15;
  assign maxi_wstrb = _sb_maxi_writedata_m_value_14;
  assign maxi_wlast = _sb_maxi_writedata_m_value_13;
  assign maxi_wvalid = _sb_maxi_writedata_valid_7;
  assign maxi_bready = 1;
  assign maxi_arsize = 2;
  assign maxi_arburst = 1;
  assign maxi_arlock = 0;
  assign maxi_arcache = 3;
  assign maxi_arprot = 0;
  assign maxi_arqos = 0;
  assign maxi_aruser = 0;
  wire [32-1:0] _maxi_rdata_sb_0;
  wire _maxi_rlast_sb_0;
  wire _maxi_rvalid_sb_0;
  wire _maxi_rready_sb_0;
  wire _sb_maxi_readdata_s_value_16;
  assign _sb_maxi_readdata_s_value_16 = maxi_rlast;
  wire [32-1:0] _sb_maxi_readdata_s_value_17;
  assign _sb_maxi_readdata_s_value_17 = maxi_rdata;
  wire [33-1:0] _sb_maxi_readdata_s_data_18;
  assign _sb_maxi_readdata_s_data_18 = { _sb_maxi_readdata_s_value_16, _sb_maxi_readdata_s_value_17 };
  wire _sb_maxi_readdata_s_valid_19;
  assign _sb_maxi_readdata_s_valid_19 = maxi_rvalid;
  wire _sb_maxi_readdata_m_ready_20;
  assign _sb_maxi_readdata_m_ready_20 = _maxi_rready_sb_0;
  reg [33-1:0] _sb_maxi_readdata_data_21;
  reg _sb_maxi_readdata_valid_22;
  wire _sb_maxi_readdata_ready_23;
  reg [33-1:0] _sb_maxi_readdata_tmp_data_24;
  reg _sb_maxi_readdata_tmp_valid_25;
  wire [33-1:0] _sb_maxi_readdata_next_data_26;
  wire _sb_maxi_readdata_next_valid_27;
  assign _sb_maxi_readdata_ready_23 = !_sb_maxi_readdata_tmp_valid_25;
  assign _sb_maxi_readdata_next_data_26 = (_sb_maxi_readdata_tmp_valid_25)? _sb_maxi_readdata_tmp_data_24 : _sb_maxi_readdata_s_data_18;
  assign _sb_maxi_readdata_next_valid_27 = _sb_maxi_readdata_tmp_valid_25 || _sb_maxi_readdata_s_valid_19;
  wire _sb_maxi_readdata_m_value_28;
  assign _sb_maxi_readdata_m_value_28 = _sb_maxi_readdata_data_21[32:32];
  wire [32-1:0] _sb_maxi_readdata_m_value_29;
  assign _sb_maxi_readdata_m_value_29 = _sb_maxi_readdata_data_21[31:0];
  assign _maxi_rdata_sb_0 = _sb_maxi_readdata_m_value_29;
  assign _maxi_rlast_sb_0 = _sb_maxi_readdata_m_value_28;
  assign _maxi_rvalid_sb_0 = _sb_maxi_readdata_valid_22;
  assign maxi_rready = _sb_maxi_readdata_ready_23;
  reg [3-1:0] _maxi_outstanding_wcount;
  wire _maxi_has_outstanding_write;
  assign _maxi_has_outstanding_write = (_maxi_outstanding_wcount > 0) || maxi_awvalid;
  reg _maxi_read_start;
  reg [8-1:0] _maxi_read_op_sel;
  reg [32-1:0] _maxi_read_global_addr;
  reg [33-1:0] _maxi_read_global_size;
  reg [32-1:0] _maxi_read_local_addr;
  reg [32-1:0] _maxi_read_local_stride;
  reg [33-1:0] _maxi_read_local_size;
  reg [32-1:0] _maxi_read_local_blocksize;
  wire _maxi_read_req_fifo_enq;
  wire [137-1:0] _maxi_read_req_fifo_wdata;
  wire _maxi_read_req_fifo_full;
  wire _maxi_read_req_fifo_almost_full;
  wire _maxi_read_req_fifo_deq;
  wire [137-1:0] _maxi_read_req_fifo_rdata;
  wire _maxi_read_req_fifo_empty;
  wire _maxi_read_req_fifo_almost_empty;

  _maxi_read_req_fifo
  inst__maxi_read_req_fifo
  (
    .CLK(CLK),
    .RST(RESETN_inv_buf),
    ._maxi_read_req_fifo_enq(_maxi_read_req_fifo_enq),
    ._maxi_read_req_fifo_wdata(_maxi_read_req_fifo_wdata),
    ._maxi_read_req_fifo_full(_maxi_read_req_fifo_full),
    ._maxi_read_req_fifo_almost_full(_maxi_read_req_fifo_almost_full),
    ._maxi_read_req_fifo_deq(_maxi_read_req_fifo_deq),
    ._maxi_read_req_fifo_rdata(_maxi_read_req_fifo_rdata),
    ._maxi_read_req_fifo_empty(_maxi_read_req_fifo_empty),
    ._maxi_read_req_fifo_almost_empty(_maxi_read_req_fifo_almost_empty)
  );

  reg [4-1:0] count__maxi_read_req_fifo;
  wire [8-1:0] _maxi_read_op_sel_fifo;
  wire [32-1:0] _maxi_read_local_addr_fifo;
  wire [32-1:0] _maxi_read_local_stride_fifo;
  wire [33-1:0] _maxi_read_local_size_fifo;
  wire [32-1:0] _maxi_read_local_blocksize_fifo;
  wire [8-1:0] unpack_read_req_op_sel_30;
  wire [32-1:0] unpack_read_req_local_addr_31;
  wire [32-1:0] unpack_read_req_local_stride_32;
  wire [33-1:0] unpack_read_req_local_size_33;
  wire [32-1:0] unpack_read_req_local_blocksize_34;
  assign unpack_read_req_op_sel_30 = _maxi_read_req_fifo_rdata[136:129];
  assign unpack_read_req_local_addr_31 = _maxi_read_req_fifo_rdata[128:97];
  assign unpack_read_req_local_stride_32 = _maxi_read_req_fifo_rdata[96:65];
  assign unpack_read_req_local_size_33 = _maxi_read_req_fifo_rdata[64:32];
  assign unpack_read_req_local_blocksize_34 = _maxi_read_req_fifo_rdata[31:0];
  assign _maxi_read_op_sel_fifo = unpack_read_req_op_sel_30;
  assign _maxi_read_local_addr_fifo = unpack_read_req_local_addr_31;
  assign _maxi_read_local_stride_fifo = unpack_read_req_local_stride_32;
  assign _maxi_read_local_size_fifo = unpack_read_req_local_size_33;
  assign _maxi_read_local_blocksize_fifo = unpack_read_req_local_blocksize_34;
  reg [8-1:0] _maxi_read_op_sel_buf;
  reg [32-1:0] _maxi_read_local_addr_buf;
  reg [32-1:0] _maxi_read_local_stride_buf;
  reg [33-1:0] _maxi_read_local_size_buf;
  reg [32-1:0] _maxi_read_local_blocksize_buf;
  reg _maxi_read_req_busy;
  reg _maxi_read_data_busy;
  wire _maxi_read_req_idle;
  wire _maxi_read_data_idle;
  wire _maxi_read_idle;
  assign _maxi_read_req_idle = !_maxi_read_start && !_maxi_read_req_busy;
  assign _maxi_read_data_idle = _maxi_read_req_fifo_empty && !_maxi_read_data_busy;
  assign _maxi_read_idle = _maxi_read_req_idle && _maxi_read_data_idle;
  reg _maxi_write_start;
  reg [8-1:0] _maxi_write_op_sel;
  reg [32-1:0] _maxi_write_global_addr;
  reg [33-1:0] _maxi_write_global_size;
  reg [32-1:0] _maxi_write_local_addr;
  reg [32-1:0] _maxi_write_local_stride;
  reg [33-1:0] _maxi_write_local_size;
  reg [32-1:0] _maxi_write_local_blocksize;
  wire _maxi_write_req_fifo_enq;
  wire [137-1:0] _maxi_write_req_fifo_wdata;
  wire _maxi_write_req_fifo_full;
  wire _maxi_write_req_fifo_almost_full;
  wire _maxi_write_req_fifo_deq;
  wire [137-1:0] _maxi_write_req_fifo_rdata;
  wire _maxi_write_req_fifo_empty;
  wire _maxi_write_req_fifo_almost_empty;

  _maxi_write_req_fifo
  inst__maxi_write_req_fifo
  (
    .CLK(CLK),
    .RST(RESETN_inv_buf),
    ._maxi_write_req_fifo_enq(_maxi_write_req_fifo_enq),
    ._maxi_write_req_fifo_wdata(_maxi_write_req_fifo_wdata),
    ._maxi_write_req_fifo_full(_maxi_write_req_fifo_full),
    ._maxi_write_req_fifo_almost_full(_maxi_write_req_fifo_almost_full),
    ._maxi_write_req_fifo_deq(_maxi_write_req_fifo_deq),
    ._maxi_write_req_fifo_rdata(_maxi_write_req_fifo_rdata),
    ._maxi_write_req_fifo_empty(_maxi_write_req_fifo_empty),
    ._maxi_write_req_fifo_almost_empty(_maxi_write_req_fifo_almost_empty)
  );

  reg [4-1:0] count__maxi_write_req_fifo;
  wire [8-1:0] _maxi_write_op_sel_fifo;
  wire [32-1:0] _maxi_write_local_addr_fifo;
  wire [32-1:0] _maxi_write_local_stride_fifo;
  wire [33-1:0] _maxi_write_size_fifo;
  wire [32-1:0] _maxi_write_local_blocksize_fifo;
  wire [8-1:0] unpack_write_req_op_sel_35;
  wire [32-1:0] unpack_write_req_local_addr_36;
  wire [32-1:0] unpack_write_req_local_stride_37;
  wire [33-1:0] unpack_write_req_size_38;
  wire [32-1:0] unpack_write_req_local_blocksize_39;
  assign unpack_write_req_op_sel_35 = _maxi_write_req_fifo_rdata[136:129];
  assign unpack_write_req_local_addr_36 = _maxi_write_req_fifo_rdata[128:97];
  assign unpack_write_req_local_stride_37 = _maxi_write_req_fifo_rdata[96:65];
  assign unpack_write_req_size_38 = _maxi_write_req_fifo_rdata[64:32];
  assign unpack_write_req_local_blocksize_39 = _maxi_write_req_fifo_rdata[31:0];
  assign _maxi_write_op_sel_fifo = unpack_write_req_op_sel_35;
  assign _maxi_write_local_addr_fifo = unpack_write_req_local_addr_36;
  assign _maxi_write_local_stride_fifo = unpack_write_req_local_stride_37;
  assign _maxi_write_size_fifo = unpack_write_req_size_38;
  assign _maxi_write_local_blocksize_fifo = unpack_write_req_local_blocksize_39;
  reg [8-1:0] _maxi_write_op_sel_buf;
  reg [32-1:0] _maxi_write_local_addr_buf;
  reg [32-1:0] _maxi_write_local_stride_buf;
  reg [33-1:0] _maxi_write_size_buf;
  reg [32-1:0] _maxi_write_local_blocksize_buf;
  reg _maxi_write_req_busy;
  reg _maxi_write_data_busy;
  wire _maxi_write_req_idle;
  wire _maxi_write_data_idle;
  wire _maxi_write_idle;
  assign _maxi_write_req_idle = !_maxi_write_start && !_maxi_write_req_busy;
  assign _maxi_write_data_idle = _maxi_write_req_fifo_empty && !_maxi_write_data_busy;
  assign _maxi_write_idle = _maxi_write_req_idle && _maxi_write_data_idle;
  reg [32-1:0] _maxi_global_base_addr;
  assign saxi_bresp = 0;
  assign saxi_rresp = 0;
  reg signed [32-1:0] _saxi_register_0;
  reg signed [32-1:0] _saxi_register_1;
  reg signed [32-1:0] _saxi_register_2;
  reg signed [32-1:0] _saxi_register_3;
  reg signed [32-1:0] _saxi_register_4;
  reg signed [32-1:0] _saxi_register_5;
  reg signed [32-1:0] _saxi_register_6;
  reg signed [32-1:0] _saxi_register_7;
  reg signed [32-1:0] _saxi_register_8;
  reg signed [32-1:0] _saxi_register_9;
  reg signed [32-1:0] _saxi_register_10;
  reg signed [32-1:0] _saxi_register_11;
  reg signed [32-1:0] _saxi_register_12;
  reg signed [32-1:0] _saxi_register_13;
  reg signed [32-1:0] _saxi_register_14;
  reg signed [32-1:0] _saxi_register_15;
  reg signed [32-1:0] _saxi_register_16;
  reg signed [32-1:0] _saxi_register_17;
  reg signed [32-1:0] _saxi_register_18;
  reg signed [32-1:0] _saxi_register_19;
  reg signed [32-1:0] _saxi_register_20;
  reg signed [32-1:0] _saxi_register_21;
  reg signed [32-1:0] _saxi_register_22;
  reg signed [32-1:0] _saxi_register_23;
  reg signed [32-1:0] _saxi_register_24;
  reg signed [32-1:0] _saxi_register_25;
  reg signed [32-1:0] _saxi_register_26;
  reg signed [32-1:0] _saxi_register_27;
  reg signed [32-1:0] _saxi_register_28;
  reg signed [32-1:0] _saxi_register_29;
  reg signed [32-1:0] _saxi_register_30;
  reg signed [32-1:0] _saxi_register_31;
  reg signed [32-1:0] _saxi_register_32;
  reg signed [32-1:0] _saxi_register_33;
  reg signed [32-1:0] _saxi_register_34;
  reg signed [32-1:0] _saxi_register_35;
  reg signed [32-1:0] _saxi_register_36;
  reg _saxi_flag_0;
  reg _saxi_flag_1;
  reg _saxi_flag_2;
  reg _saxi_flag_3;
  reg _saxi_flag_4;
  reg _saxi_flag_5;
  reg _saxi_flag_6;
  reg _saxi_flag_7;
  reg _saxi_flag_8;
  reg _saxi_flag_9;
  reg _saxi_flag_10;
  reg _saxi_flag_11;
  reg _saxi_flag_12;
  reg _saxi_flag_13;
  reg _saxi_flag_14;
  reg _saxi_flag_15;
  reg _saxi_flag_16;
  reg _saxi_flag_17;
  reg _saxi_flag_18;
  reg _saxi_flag_19;
  reg _saxi_flag_20;
  reg _saxi_flag_21;
  reg _saxi_flag_22;
  reg _saxi_flag_23;
  reg _saxi_flag_24;
  reg _saxi_flag_25;
  reg _saxi_flag_26;
  reg _saxi_flag_27;
  reg _saxi_flag_28;
  reg _saxi_flag_29;
  reg _saxi_flag_30;
  reg _saxi_flag_31;
  reg _saxi_flag_32;
  reg _saxi_flag_33;
  reg _saxi_flag_34;
  reg _saxi_flag_35;
  reg _saxi_flag_36;
  reg signed [32-1:0] _saxi_resetval_0;
  reg signed [32-1:0] _saxi_resetval_1;
  reg signed [32-1:0] _saxi_resetval_2;
  reg signed [32-1:0] _saxi_resetval_3;
  reg signed [32-1:0] _saxi_resetval_4;
  reg signed [32-1:0] _saxi_resetval_5;
  reg signed [32-1:0] _saxi_resetval_6;
  reg signed [32-1:0] _saxi_resetval_7;
  reg signed [32-1:0] _saxi_resetval_8;
  reg signed [32-1:0] _saxi_resetval_9;
  reg signed [32-1:0] _saxi_resetval_10;
  reg signed [32-1:0] _saxi_resetval_11;
  reg signed [32-1:0] _saxi_resetval_12;
  reg signed [32-1:0] _saxi_resetval_13;
  reg signed [32-1:0] _saxi_resetval_14;
  reg signed [32-1:0] _saxi_resetval_15;
  reg signed [32-1:0] _saxi_resetval_16;
  reg signed [32-1:0] _saxi_resetval_17;
  reg signed [32-1:0] _saxi_resetval_18;
  reg signed [32-1:0] _saxi_resetval_19;
  reg signed [32-1:0] _saxi_resetval_20;
  reg signed [32-1:0] _saxi_resetval_21;
  reg signed [32-1:0] _saxi_resetval_22;
  reg signed [32-1:0] _saxi_resetval_23;
  reg signed [32-1:0] _saxi_resetval_24;
  reg signed [32-1:0] _saxi_resetval_25;
  reg signed [32-1:0] _saxi_resetval_26;
  reg signed [32-1:0] _saxi_resetval_27;
  reg signed [32-1:0] _saxi_resetval_28;
  reg signed [32-1:0] _saxi_resetval_29;
  reg signed [32-1:0] _saxi_resetval_30;
  reg signed [32-1:0] _saxi_resetval_31;
  reg signed [32-1:0] _saxi_resetval_32;
  reg signed [32-1:0] _saxi_resetval_33;
  reg signed [32-1:0] _saxi_resetval_34;
  reg signed [32-1:0] _saxi_resetval_35;
  reg signed [32-1:0] _saxi_resetval_36;
  localparam _saxi_maskwidth = 6;
  localparam _saxi_mask = { _saxi_maskwidth{ 1'd1 } };
  localparam _saxi_shift = 2;
  reg [32-1:0] _saxi_register_fsm;
  localparam _saxi_register_fsm_init = 0;
  reg [32-1:0] addr_40;
  reg writevalid_41;
  reg readvalid_42;
  reg prev_awvalid_43;
  reg prev_arvalid_44;
  assign saxi_awready = (_saxi_register_fsm == 0) && (!writevalid_41 && !readvalid_42 && !saxi_bvalid && prev_awvalid_43);
  assign saxi_arready = (_saxi_register_fsm == 0) && (!readvalid_42 && !writevalid_41 && prev_arvalid_44 && !prev_awvalid_43);
  reg [_saxi_maskwidth-1:0] axis_maskaddr_45;
  wire signed [32-1:0] axislite_rdata_46;
  assign axislite_rdata_46 = (axis_maskaddr_45 == 0)? _saxi_register_0 : 
                             (axis_maskaddr_45 == 1)? _saxi_register_1 : 
                             (axis_maskaddr_45 == 2)? _saxi_register_2 : 
                             (axis_maskaddr_45 == 3)? _saxi_register_3 : 
                             (axis_maskaddr_45 == 4)? _saxi_register_4 : 
                             (axis_maskaddr_45 == 5)? _saxi_register_5 : 
                             (axis_maskaddr_45 == 6)? _saxi_register_6 : 
                             (axis_maskaddr_45 == 7)? _saxi_register_7 : 
                             (axis_maskaddr_45 == 8)? _saxi_register_8 : 
                             (axis_maskaddr_45 == 9)? _saxi_register_9 : 
                             (axis_maskaddr_45 == 10)? _saxi_register_10 : 
                             (axis_maskaddr_45 == 11)? _saxi_register_11 : 
                             (axis_maskaddr_45 == 12)? _saxi_register_12 : 
                             (axis_maskaddr_45 == 13)? _saxi_register_13 : 
                             (axis_maskaddr_45 == 14)? _saxi_register_14 : 
                             (axis_maskaddr_45 == 15)? _saxi_register_15 : 
                             (axis_maskaddr_45 == 16)? _saxi_register_16 : 
                             (axis_maskaddr_45 == 17)? _saxi_register_17 : 
                             (axis_maskaddr_45 == 18)? _saxi_register_18 : 
                             (axis_maskaddr_45 == 19)? _saxi_register_19 : 
                             (axis_maskaddr_45 == 20)? _saxi_register_20 : 
                             (axis_maskaddr_45 == 21)? _saxi_register_21 : 
                             (axis_maskaddr_45 == 22)? _saxi_register_22 : 
                             (axis_maskaddr_45 == 23)? _saxi_register_23 : 
                             (axis_maskaddr_45 == 24)? _saxi_register_24 : 
                             (axis_maskaddr_45 == 25)? _saxi_register_25 : 
                             (axis_maskaddr_45 == 26)? _saxi_register_26 : 
                             (axis_maskaddr_45 == 27)? _saxi_register_27 : 
                             (axis_maskaddr_45 == 28)? _saxi_register_28 : 
                             (axis_maskaddr_45 == 29)? _saxi_register_29 : 
                             (axis_maskaddr_45 == 30)? _saxi_register_30 : 
                             (axis_maskaddr_45 == 31)? _saxi_register_31 : 
                             (axis_maskaddr_45 == 32)? _saxi_register_32 : 
                             (axis_maskaddr_45 == 33)? _saxi_register_33 : 
                             (axis_maskaddr_45 == 34)? _saxi_register_34 : 
                             (axis_maskaddr_45 == 35)? _saxi_register_35 : 
                             (axis_maskaddr_45 == 36)? _saxi_register_36 : 'hx;
  wire axislite_flag_47;
  assign axislite_flag_47 = (axis_maskaddr_45 == 0)? _saxi_flag_0 : 
                            (axis_maskaddr_45 == 1)? _saxi_flag_1 : 
                            (axis_maskaddr_45 == 2)? _saxi_flag_2 : 
                            (axis_maskaddr_45 == 3)? _saxi_flag_3 : 
                            (axis_maskaddr_45 == 4)? _saxi_flag_4 : 
                            (axis_maskaddr_45 == 5)? _saxi_flag_5 : 
                            (axis_maskaddr_45 == 6)? _saxi_flag_6 : 
                            (axis_maskaddr_45 == 7)? _saxi_flag_7 : 
                            (axis_maskaddr_45 == 8)? _saxi_flag_8 : 
                            (axis_maskaddr_45 == 9)? _saxi_flag_9 : 
                            (axis_maskaddr_45 == 10)? _saxi_flag_10 : 
                            (axis_maskaddr_45 == 11)? _saxi_flag_11 : 
                            (axis_maskaddr_45 == 12)? _saxi_flag_12 : 
                            (axis_maskaddr_45 == 13)? _saxi_flag_13 : 
                            (axis_maskaddr_45 == 14)? _saxi_flag_14 : 
                            (axis_maskaddr_45 == 15)? _saxi_flag_15 : 
                            (axis_maskaddr_45 == 16)? _saxi_flag_16 : 
                            (axis_maskaddr_45 == 17)? _saxi_flag_17 : 
                            (axis_maskaddr_45 == 18)? _saxi_flag_18 : 
                            (axis_maskaddr_45 == 19)? _saxi_flag_19 : 
                            (axis_maskaddr_45 == 20)? _saxi_flag_20 : 
                            (axis_maskaddr_45 == 21)? _saxi_flag_21 : 
                            (axis_maskaddr_45 == 22)? _saxi_flag_22 : 
                            (axis_maskaddr_45 == 23)? _saxi_flag_23 : 
                            (axis_maskaddr_45 == 24)? _saxi_flag_24 : 
                            (axis_maskaddr_45 == 25)? _saxi_flag_25 : 
                            (axis_maskaddr_45 == 26)? _saxi_flag_26 : 
                            (axis_maskaddr_45 == 27)? _saxi_flag_27 : 
                            (axis_maskaddr_45 == 28)? _saxi_flag_28 : 
                            (axis_maskaddr_45 == 29)? _saxi_flag_29 : 
                            (axis_maskaddr_45 == 30)? _saxi_flag_30 : 
                            (axis_maskaddr_45 == 31)? _saxi_flag_31 : 
                            (axis_maskaddr_45 == 32)? _saxi_flag_32 : 
                            (axis_maskaddr_45 == 33)? _saxi_flag_33 : 
                            (axis_maskaddr_45 == 34)? _saxi_flag_34 : 
                            (axis_maskaddr_45 == 35)? _saxi_flag_35 : 
                            (axis_maskaddr_45 == 36)? _saxi_flag_36 : 'hx;
  wire signed [32-1:0] axislite_resetval_48;
  assign axislite_resetval_48 = (axis_maskaddr_45 == 0)? _saxi_resetval_0 : 
                                (axis_maskaddr_45 == 1)? _saxi_resetval_1 : 
                                (axis_maskaddr_45 == 2)? _saxi_resetval_2 : 
                                (axis_maskaddr_45 == 3)? _saxi_resetval_3 : 
                                (axis_maskaddr_45 == 4)? _saxi_resetval_4 : 
                                (axis_maskaddr_45 == 5)? _saxi_resetval_5 : 
                                (axis_maskaddr_45 == 6)? _saxi_resetval_6 : 
                                (axis_maskaddr_45 == 7)? _saxi_resetval_7 : 
                                (axis_maskaddr_45 == 8)? _saxi_resetval_8 : 
                                (axis_maskaddr_45 == 9)? _saxi_resetval_9 : 
                                (axis_maskaddr_45 == 10)? _saxi_resetval_10 : 
                                (axis_maskaddr_45 == 11)? _saxi_resetval_11 : 
                                (axis_maskaddr_45 == 12)? _saxi_resetval_12 : 
                                (axis_maskaddr_45 == 13)? _saxi_resetval_13 : 
                                (axis_maskaddr_45 == 14)? _saxi_resetval_14 : 
                                (axis_maskaddr_45 == 15)? _saxi_resetval_15 : 
                                (axis_maskaddr_45 == 16)? _saxi_resetval_16 : 
                                (axis_maskaddr_45 == 17)? _saxi_resetval_17 : 
                                (axis_maskaddr_45 == 18)? _saxi_resetval_18 : 
                                (axis_maskaddr_45 == 19)? _saxi_resetval_19 : 
                                (axis_maskaddr_45 == 20)? _saxi_resetval_20 : 
                                (axis_maskaddr_45 == 21)? _saxi_resetval_21 : 
                                (axis_maskaddr_45 == 22)? _saxi_resetval_22 : 
                                (axis_maskaddr_45 == 23)? _saxi_resetval_23 : 
                                (axis_maskaddr_45 == 24)? _saxi_resetval_24 : 
                                (axis_maskaddr_45 == 25)? _saxi_resetval_25 : 
                                (axis_maskaddr_45 == 26)? _saxi_resetval_26 : 
                                (axis_maskaddr_45 == 27)? _saxi_resetval_27 : 
                                (axis_maskaddr_45 == 28)? _saxi_resetval_28 : 
                                (axis_maskaddr_45 == 29)? _saxi_resetval_29 : 
                                (axis_maskaddr_45 == 30)? _saxi_resetval_30 : 
                                (axis_maskaddr_45 == 31)? _saxi_resetval_31 : 
                                (axis_maskaddr_45 == 32)? _saxi_resetval_32 : 
                                (axis_maskaddr_45 == 33)? _saxi_resetval_33 : 
                                (axis_maskaddr_45 == 34)? _saxi_resetval_34 : 
                                (axis_maskaddr_45 == 35)? _saxi_resetval_35 : 
                                (axis_maskaddr_45 == 36)? _saxi_resetval_36 : 'hx;
  reg _saxi_rdata_cond_0_1;
  assign saxi_wready = _saxi_register_fsm == 3;
  wire maxi_idle;
  assign maxi_idle = _maxi_write_idle & _maxi_read_idle;
  wire sw_rst_logic;
  assign sw_rst_logic = maxi_idle & _saxi_register_6;
  wire rst_logic;
  assign rst_logic = RESETN_inv_buf | sw_rst_logic;
  reg RST;
  reg _rst_logic_1;
  reg _rst_logic_2;
  wire signed [32-1:0] irq_49;
  assign irq_49 = _saxi_register_9 & _saxi_register_10;
  wire irq_busy;
  assign irq_busy = _saxi_register_5[0];
  reg irq_busy_edge_50;
  wire irq_busy_edge_51;
  assign irq_busy_edge_51 = irq_busy_edge_50 & !irq_busy;
  wire irq_extern;
  assign irq_extern = |_saxi_register_7;
  reg irq_extern_edge_52;
  wire irq_extern_edge_53;
  assign irq_extern_edge_53 = !irq_extern_edge_52 & irq_extern;
  wire [14-1:0] ram_w16_l32768_id0_0_0_addr;
  wire [16-1:0] ram_w16_l32768_id0_0_0_rdata;
  wire [16-1:0] ram_w16_l32768_id0_0_0_wdata;
  wire ram_w16_l32768_id0_0_0_wenable;
  wire ram_w16_l32768_id0_0_0_enable;
  wire [14-1:0] ram_w16_l32768_id0_0_1_addr;
  wire [16-1:0] ram_w16_l32768_id0_0_1_rdata;
  wire [16-1:0] ram_w16_l32768_id0_0_1_wdata;
  wire ram_w16_l32768_id0_0_1_wenable;
  wire ram_w16_l32768_id0_0_1_enable;
  assign ram_w16_l32768_id0_0_0_wdata = 'hx;
  assign ram_w16_l32768_id0_0_0_wenable = 0;

  ram_w16_l32768_id0_0
  inst_ram_w16_l32768_id0_0
  (
    .CLK(CLK),
    .ram_w16_l32768_id0_0_0_addr(ram_w16_l32768_id0_0_0_addr),
    .ram_w16_l32768_id0_0_0_rdata(ram_w16_l32768_id0_0_0_rdata),
    .ram_w16_l32768_id0_0_0_wdata(ram_w16_l32768_id0_0_0_wdata),
    .ram_w16_l32768_id0_0_0_wenable(ram_w16_l32768_id0_0_0_wenable),
    .ram_w16_l32768_id0_0_0_enable(ram_w16_l32768_id0_0_0_enable),
    .ram_w16_l32768_id0_0_1_addr(ram_w16_l32768_id0_0_1_addr),
    .ram_w16_l32768_id0_0_1_rdata(ram_w16_l32768_id0_0_1_rdata),
    .ram_w16_l32768_id0_0_1_wdata(ram_w16_l32768_id0_0_1_wdata),
    .ram_w16_l32768_id0_0_1_wenable(ram_w16_l32768_id0_0_1_wenable),
    .ram_w16_l32768_id0_0_1_enable(ram_w16_l32768_id0_0_1_enable)
  );

  wire [14-1:0] ram_w16_l32768_id0_1_0_addr;
  wire [16-1:0] ram_w16_l32768_id0_1_0_rdata;
  wire [16-1:0] ram_w16_l32768_id0_1_0_wdata;
  wire ram_w16_l32768_id0_1_0_wenable;
  wire ram_w16_l32768_id0_1_0_enable;
  wire [14-1:0] ram_w16_l32768_id0_1_1_addr;
  wire [16-1:0] ram_w16_l32768_id0_1_1_rdata;
  wire [16-1:0] ram_w16_l32768_id0_1_1_wdata;
  wire ram_w16_l32768_id0_1_1_wenable;
  wire ram_w16_l32768_id0_1_1_enable;
  assign ram_w16_l32768_id0_1_0_wdata = 'hx;
  assign ram_w16_l32768_id0_1_0_wenable = 0;

  ram_w16_l32768_id0_1
  inst_ram_w16_l32768_id0_1
  (
    .CLK(CLK),
    .ram_w16_l32768_id0_1_0_addr(ram_w16_l32768_id0_1_0_addr),
    .ram_w16_l32768_id0_1_0_rdata(ram_w16_l32768_id0_1_0_rdata),
    .ram_w16_l32768_id0_1_0_wdata(ram_w16_l32768_id0_1_0_wdata),
    .ram_w16_l32768_id0_1_0_wenable(ram_w16_l32768_id0_1_0_wenable),
    .ram_w16_l32768_id0_1_0_enable(ram_w16_l32768_id0_1_0_enable),
    .ram_w16_l32768_id0_1_1_addr(ram_w16_l32768_id0_1_1_addr),
    .ram_w16_l32768_id0_1_1_rdata(ram_w16_l32768_id0_1_1_rdata),
    .ram_w16_l32768_id0_1_1_wdata(ram_w16_l32768_id0_1_1_wdata),
    .ram_w16_l32768_id0_1_1_wenable(ram_w16_l32768_id0_1_1_wenable),
    .ram_w16_l32768_id0_1_1_enable(ram_w16_l32768_id0_1_1_enable)
  );

  wire [12-1:0] ram_w16_l8192_id0_0_0_addr;
  wire [16-1:0] ram_w16_l8192_id0_0_0_rdata;
  wire [16-1:0] ram_w16_l8192_id0_0_0_wdata;
  wire ram_w16_l8192_id0_0_0_wenable;
  wire ram_w16_l8192_id0_0_0_enable;
  wire [12-1:0] ram_w16_l8192_id0_0_1_addr;
  wire [16-1:0] ram_w16_l8192_id0_0_1_rdata;
  wire [16-1:0] ram_w16_l8192_id0_0_1_wdata;
  wire ram_w16_l8192_id0_0_1_wenable;
  wire ram_w16_l8192_id0_0_1_enable;

  ram_w16_l8192_id0_0
  inst_ram_w16_l8192_id0_0
  (
    .CLK(CLK),
    .ram_w16_l8192_id0_0_0_addr(ram_w16_l8192_id0_0_0_addr),
    .ram_w16_l8192_id0_0_0_rdata(ram_w16_l8192_id0_0_0_rdata),
    .ram_w16_l8192_id0_0_0_wdata(ram_w16_l8192_id0_0_0_wdata),
    .ram_w16_l8192_id0_0_0_wenable(ram_w16_l8192_id0_0_0_wenable),
    .ram_w16_l8192_id0_0_0_enable(ram_w16_l8192_id0_0_0_enable),
    .ram_w16_l8192_id0_0_1_addr(ram_w16_l8192_id0_0_1_addr),
    .ram_w16_l8192_id0_0_1_rdata(ram_w16_l8192_id0_0_1_rdata),
    .ram_w16_l8192_id0_0_1_wdata(ram_w16_l8192_id0_0_1_wdata),
    .ram_w16_l8192_id0_0_1_wenable(ram_w16_l8192_id0_0_1_wenable),
    .ram_w16_l8192_id0_0_1_enable(ram_w16_l8192_id0_0_1_enable)
  );

  wire [12-1:0] ram_w16_l8192_id0_1_0_addr;
  wire [16-1:0] ram_w16_l8192_id0_1_0_rdata;
  wire [16-1:0] ram_w16_l8192_id0_1_0_wdata;
  wire ram_w16_l8192_id0_1_0_wenable;
  wire ram_w16_l8192_id0_1_0_enable;
  wire [12-1:0] ram_w16_l8192_id0_1_1_addr;
  wire [16-1:0] ram_w16_l8192_id0_1_1_rdata;
  wire [16-1:0] ram_w16_l8192_id0_1_1_wdata;
  wire ram_w16_l8192_id0_1_1_wenable;
  wire ram_w16_l8192_id0_1_1_enable;

  ram_w16_l8192_id0_1
  inst_ram_w16_l8192_id0_1
  (
    .CLK(CLK),
    .ram_w16_l8192_id0_1_0_addr(ram_w16_l8192_id0_1_0_addr),
    .ram_w16_l8192_id0_1_0_rdata(ram_w16_l8192_id0_1_0_rdata),
    .ram_w16_l8192_id0_1_0_wdata(ram_w16_l8192_id0_1_0_wdata),
    .ram_w16_l8192_id0_1_0_wenable(ram_w16_l8192_id0_1_0_wenable),
    .ram_w16_l8192_id0_1_0_enable(ram_w16_l8192_id0_1_0_enable),
    .ram_w16_l8192_id0_1_1_addr(ram_w16_l8192_id0_1_1_addr),
    .ram_w16_l8192_id0_1_1_rdata(ram_w16_l8192_id0_1_1_rdata),
    .ram_w16_l8192_id0_1_1_wdata(ram_w16_l8192_id0_1_1_wdata),
    .ram_w16_l8192_id0_1_1_wenable(ram_w16_l8192_id0_1_1_wenable),
    .ram_w16_l8192_id0_1_1_enable(ram_w16_l8192_id0_1_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id0_0_0_addr;
  wire [16-1:0] ram_w16_l512_id0_0_0_rdata;
  wire [16-1:0] ram_w16_l512_id0_0_0_wdata;
  wire ram_w16_l512_id0_0_0_wenable;
  wire ram_w16_l512_id0_0_0_enable;
  wire [8-1:0] ram_w16_l512_id0_0_1_addr;
  wire [16-1:0] ram_w16_l512_id0_0_1_rdata;
  wire [16-1:0] ram_w16_l512_id0_0_1_wdata;
  wire ram_w16_l512_id0_0_1_wenable;
  wire ram_w16_l512_id0_0_1_enable;

  ram_w16_l512_id0_0
  inst_ram_w16_l512_id0_0
  (
    .CLK(CLK),
    .ram_w16_l512_id0_0_0_addr(ram_w16_l512_id0_0_0_addr),
    .ram_w16_l512_id0_0_0_rdata(ram_w16_l512_id0_0_0_rdata),
    .ram_w16_l512_id0_0_0_wdata(ram_w16_l512_id0_0_0_wdata),
    .ram_w16_l512_id0_0_0_wenable(ram_w16_l512_id0_0_0_wenable),
    .ram_w16_l512_id0_0_0_enable(ram_w16_l512_id0_0_0_enable),
    .ram_w16_l512_id0_0_1_addr(ram_w16_l512_id0_0_1_addr),
    .ram_w16_l512_id0_0_1_rdata(ram_w16_l512_id0_0_1_rdata),
    .ram_w16_l512_id0_0_1_wdata(ram_w16_l512_id0_0_1_wdata),
    .ram_w16_l512_id0_0_1_wenable(ram_w16_l512_id0_0_1_wenable),
    .ram_w16_l512_id0_0_1_enable(ram_w16_l512_id0_0_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id0_1_0_addr;
  wire [16-1:0] ram_w16_l512_id0_1_0_rdata;
  wire [16-1:0] ram_w16_l512_id0_1_0_wdata;
  wire ram_w16_l512_id0_1_0_wenable;
  wire ram_w16_l512_id0_1_0_enable;
  wire [8-1:0] ram_w16_l512_id0_1_1_addr;
  wire [16-1:0] ram_w16_l512_id0_1_1_rdata;
  wire [16-1:0] ram_w16_l512_id0_1_1_wdata;
  wire ram_w16_l512_id0_1_1_wenable;
  wire ram_w16_l512_id0_1_1_enable;

  ram_w16_l512_id0_1
  inst_ram_w16_l512_id0_1
  (
    .CLK(CLK),
    .ram_w16_l512_id0_1_0_addr(ram_w16_l512_id0_1_0_addr),
    .ram_w16_l512_id0_1_0_rdata(ram_w16_l512_id0_1_0_rdata),
    .ram_w16_l512_id0_1_0_wdata(ram_w16_l512_id0_1_0_wdata),
    .ram_w16_l512_id0_1_0_wenable(ram_w16_l512_id0_1_0_wenable),
    .ram_w16_l512_id0_1_0_enable(ram_w16_l512_id0_1_0_enable),
    .ram_w16_l512_id0_1_1_addr(ram_w16_l512_id0_1_1_addr),
    .ram_w16_l512_id0_1_1_rdata(ram_w16_l512_id0_1_1_rdata),
    .ram_w16_l512_id0_1_1_wdata(ram_w16_l512_id0_1_1_wdata),
    .ram_w16_l512_id0_1_1_wenable(ram_w16_l512_id0_1_1_wenable),
    .ram_w16_l512_id0_1_1_enable(ram_w16_l512_id0_1_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id1_0_0_addr;
  wire [16-1:0] ram_w16_l512_id1_0_0_rdata;
  wire [16-1:0] ram_w16_l512_id1_0_0_wdata;
  wire ram_w16_l512_id1_0_0_wenable;
  wire ram_w16_l512_id1_0_0_enable;
  wire [8-1:0] ram_w16_l512_id1_0_1_addr;
  wire [16-1:0] ram_w16_l512_id1_0_1_rdata;
  wire [16-1:0] ram_w16_l512_id1_0_1_wdata;
  wire ram_w16_l512_id1_0_1_wenable;
  wire ram_w16_l512_id1_0_1_enable;
  assign ram_w16_l512_id1_0_0_wdata = 'hx;
  assign ram_w16_l512_id1_0_0_wenable = 0;

  ram_w16_l512_id1_0
  inst_ram_w16_l512_id1_0
  (
    .CLK(CLK),
    .ram_w16_l512_id1_0_0_addr(ram_w16_l512_id1_0_0_addr),
    .ram_w16_l512_id1_0_0_rdata(ram_w16_l512_id1_0_0_rdata),
    .ram_w16_l512_id1_0_0_wdata(ram_w16_l512_id1_0_0_wdata),
    .ram_w16_l512_id1_0_0_wenable(ram_w16_l512_id1_0_0_wenable),
    .ram_w16_l512_id1_0_0_enable(ram_w16_l512_id1_0_0_enable),
    .ram_w16_l512_id1_0_1_addr(ram_w16_l512_id1_0_1_addr),
    .ram_w16_l512_id1_0_1_rdata(ram_w16_l512_id1_0_1_rdata),
    .ram_w16_l512_id1_0_1_wdata(ram_w16_l512_id1_0_1_wdata),
    .ram_w16_l512_id1_0_1_wenable(ram_w16_l512_id1_0_1_wenable),
    .ram_w16_l512_id1_0_1_enable(ram_w16_l512_id1_0_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id1_1_0_addr;
  wire [16-1:0] ram_w16_l512_id1_1_0_rdata;
  wire [16-1:0] ram_w16_l512_id1_1_0_wdata;
  wire ram_w16_l512_id1_1_0_wenable;
  wire ram_w16_l512_id1_1_0_enable;
  wire [8-1:0] ram_w16_l512_id1_1_1_addr;
  wire [16-1:0] ram_w16_l512_id1_1_1_rdata;
  wire [16-1:0] ram_w16_l512_id1_1_1_wdata;
  wire ram_w16_l512_id1_1_1_wenable;
  wire ram_w16_l512_id1_1_1_enable;
  assign ram_w16_l512_id1_1_0_wdata = 'hx;
  assign ram_w16_l512_id1_1_0_wenable = 0;

  ram_w16_l512_id1_1
  inst_ram_w16_l512_id1_1
  (
    .CLK(CLK),
    .ram_w16_l512_id1_1_0_addr(ram_w16_l512_id1_1_0_addr),
    .ram_w16_l512_id1_1_0_rdata(ram_w16_l512_id1_1_0_rdata),
    .ram_w16_l512_id1_1_0_wdata(ram_w16_l512_id1_1_0_wdata),
    .ram_w16_l512_id1_1_0_wenable(ram_w16_l512_id1_1_0_wenable),
    .ram_w16_l512_id1_1_0_enable(ram_w16_l512_id1_1_0_enable),
    .ram_w16_l512_id1_1_1_addr(ram_w16_l512_id1_1_1_addr),
    .ram_w16_l512_id1_1_1_rdata(ram_w16_l512_id1_1_1_rdata),
    .ram_w16_l512_id1_1_1_wdata(ram_w16_l512_id1_1_1_wdata),
    .ram_w16_l512_id1_1_1_wenable(ram_w16_l512_id1_1_1_wenable),
    .ram_w16_l512_id1_1_1_enable(ram_w16_l512_id1_1_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id2_0_0_addr;
  wire [16-1:0] ram_w16_l512_id2_0_0_rdata;
  wire [16-1:0] ram_w16_l512_id2_0_0_wdata;
  wire ram_w16_l512_id2_0_0_wenable;
  wire ram_w16_l512_id2_0_0_enable;
  wire [8-1:0] ram_w16_l512_id2_0_1_addr;
  wire [16-1:0] ram_w16_l512_id2_0_1_rdata;
  wire [16-1:0] ram_w16_l512_id2_0_1_wdata;
  wire ram_w16_l512_id2_0_1_wenable;
  wire ram_w16_l512_id2_0_1_enable;
  assign ram_w16_l512_id2_0_0_wdata = 'hx;
  assign ram_w16_l512_id2_0_0_wenable = 0;

  ram_w16_l512_id2_0
  inst_ram_w16_l512_id2_0
  (
    .CLK(CLK),
    .ram_w16_l512_id2_0_0_addr(ram_w16_l512_id2_0_0_addr),
    .ram_w16_l512_id2_0_0_rdata(ram_w16_l512_id2_0_0_rdata),
    .ram_w16_l512_id2_0_0_wdata(ram_w16_l512_id2_0_0_wdata),
    .ram_w16_l512_id2_0_0_wenable(ram_w16_l512_id2_0_0_wenable),
    .ram_w16_l512_id2_0_0_enable(ram_w16_l512_id2_0_0_enable),
    .ram_w16_l512_id2_0_1_addr(ram_w16_l512_id2_0_1_addr),
    .ram_w16_l512_id2_0_1_rdata(ram_w16_l512_id2_0_1_rdata),
    .ram_w16_l512_id2_0_1_wdata(ram_w16_l512_id2_0_1_wdata),
    .ram_w16_l512_id2_0_1_wenable(ram_w16_l512_id2_0_1_wenable),
    .ram_w16_l512_id2_0_1_enable(ram_w16_l512_id2_0_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id2_1_0_addr;
  wire [16-1:0] ram_w16_l512_id2_1_0_rdata;
  wire [16-1:0] ram_w16_l512_id2_1_0_wdata;
  wire ram_w16_l512_id2_1_0_wenable;
  wire ram_w16_l512_id2_1_0_enable;
  wire [8-1:0] ram_w16_l512_id2_1_1_addr;
  wire [16-1:0] ram_w16_l512_id2_1_1_rdata;
  wire [16-1:0] ram_w16_l512_id2_1_1_wdata;
  wire ram_w16_l512_id2_1_1_wenable;
  wire ram_w16_l512_id2_1_1_enable;
  assign ram_w16_l512_id2_1_0_wdata = 'hx;
  assign ram_w16_l512_id2_1_0_wenable = 0;

  ram_w16_l512_id2_1
  inst_ram_w16_l512_id2_1
  (
    .CLK(CLK),
    .ram_w16_l512_id2_1_0_addr(ram_w16_l512_id2_1_0_addr),
    .ram_w16_l512_id2_1_0_rdata(ram_w16_l512_id2_1_0_rdata),
    .ram_w16_l512_id2_1_0_wdata(ram_w16_l512_id2_1_0_wdata),
    .ram_w16_l512_id2_1_0_wenable(ram_w16_l512_id2_1_0_wenable),
    .ram_w16_l512_id2_1_0_enable(ram_w16_l512_id2_1_0_enable),
    .ram_w16_l512_id2_1_1_addr(ram_w16_l512_id2_1_1_addr),
    .ram_w16_l512_id2_1_1_rdata(ram_w16_l512_id2_1_1_rdata),
    .ram_w16_l512_id2_1_1_wdata(ram_w16_l512_id2_1_1_wdata),
    .ram_w16_l512_id2_1_1_wenable(ram_w16_l512_id2_1_1_wenable),
    .ram_w16_l512_id2_1_1_enable(ram_w16_l512_id2_1_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id3_0_0_addr;
  wire [16-1:0] ram_w16_l512_id3_0_0_rdata;
  wire [16-1:0] ram_w16_l512_id3_0_0_wdata;
  wire ram_w16_l512_id3_0_0_wenable;
  wire ram_w16_l512_id3_0_0_enable;
  wire [8-1:0] ram_w16_l512_id3_0_1_addr;
  wire [16-1:0] ram_w16_l512_id3_0_1_rdata;
  wire [16-1:0] ram_w16_l512_id3_0_1_wdata;
  wire ram_w16_l512_id3_0_1_wenable;
  wire ram_w16_l512_id3_0_1_enable;
  assign ram_w16_l512_id3_0_0_wdata = 'hx;
  assign ram_w16_l512_id3_0_0_wenable = 0;

  ram_w16_l512_id3_0
  inst_ram_w16_l512_id3_0
  (
    .CLK(CLK),
    .ram_w16_l512_id3_0_0_addr(ram_w16_l512_id3_0_0_addr),
    .ram_w16_l512_id3_0_0_rdata(ram_w16_l512_id3_0_0_rdata),
    .ram_w16_l512_id3_0_0_wdata(ram_w16_l512_id3_0_0_wdata),
    .ram_w16_l512_id3_0_0_wenable(ram_w16_l512_id3_0_0_wenable),
    .ram_w16_l512_id3_0_0_enable(ram_w16_l512_id3_0_0_enable),
    .ram_w16_l512_id3_0_1_addr(ram_w16_l512_id3_0_1_addr),
    .ram_w16_l512_id3_0_1_rdata(ram_w16_l512_id3_0_1_rdata),
    .ram_w16_l512_id3_0_1_wdata(ram_w16_l512_id3_0_1_wdata),
    .ram_w16_l512_id3_0_1_wenable(ram_w16_l512_id3_0_1_wenable),
    .ram_w16_l512_id3_0_1_enable(ram_w16_l512_id3_0_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id3_1_0_addr;
  wire [16-1:0] ram_w16_l512_id3_1_0_rdata;
  wire [16-1:0] ram_w16_l512_id3_1_0_wdata;
  wire ram_w16_l512_id3_1_0_wenable;
  wire ram_w16_l512_id3_1_0_enable;
  wire [8-1:0] ram_w16_l512_id3_1_1_addr;
  wire [16-1:0] ram_w16_l512_id3_1_1_rdata;
  wire [16-1:0] ram_w16_l512_id3_1_1_wdata;
  wire ram_w16_l512_id3_1_1_wenable;
  wire ram_w16_l512_id3_1_1_enable;
  assign ram_w16_l512_id3_1_0_wdata = 'hx;
  assign ram_w16_l512_id3_1_0_wenable = 0;

  ram_w16_l512_id3_1
  inst_ram_w16_l512_id3_1
  (
    .CLK(CLK),
    .ram_w16_l512_id3_1_0_addr(ram_w16_l512_id3_1_0_addr),
    .ram_w16_l512_id3_1_0_rdata(ram_w16_l512_id3_1_0_rdata),
    .ram_w16_l512_id3_1_0_wdata(ram_w16_l512_id3_1_0_wdata),
    .ram_w16_l512_id3_1_0_wenable(ram_w16_l512_id3_1_0_wenable),
    .ram_w16_l512_id3_1_0_enable(ram_w16_l512_id3_1_0_enable),
    .ram_w16_l512_id3_1_1_addr(ram_w16_l512_id3_1_1_addr),
    .ram_w16_l512_id3_1_1_rdata(ram_w16_l512_id3_1_1_rdata),
    .ram_w16_l512_id3_1_1_wdata(ram_w16_l512_id3_1_1_wdata),
    .ram_w16_l512_id3_1_1_wenable(ram_w16_l512_id3_1_1_wenable),
    .ram_w16_l512_id3_1_1_enable(ram_w16_l512_id3_1_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id4_0_0_addr;
  wire [16-1:0] ram_w16_l512_id4_0_0_rdata;
  wire [16-1:0] ram_w16_l512_id4_0_0_wdata;
  wire ram_w16_l512_id4_0_0_wenable;
  wire ram_w16_l512_id4_0_0_enable;
  wire [8-1:0] ram_w16_l512_id4_0_1_addr;
  wire [16-1:0] ram_w16_l512_id4_0_1_rdata;
  wire [16-1:0] ram_w16_l512_id4_0_1_wdata;
  wire ram_w16_l512_id4_0_1_wenable;
  wire ram_w16_l512_id4_0_1_enable;
  assign ram_w16_l512_id4_0_0_wdata = 'hx;
  assign ram_w16_l512_id4_0_0_wenable = 0;

  ram_w16_l512_id4_0
  inst_ram_w16_l512_id4_0
  (
    .CLK(CLK),
    .ram_w16_l512_id4_0_0_addr(ram_w16_l512_id4_0_0_addr),
    .ram_w16_l512_id4_0_0_rdata(ram_w16_l512_id4_0_0_rdata),
    .ram_w16_l512_id4_0_0_wdata(ram_w16_l512_id4_0_0_wdata),
    .ram_w16_l512_id4_0_0_wenable(ram_w16_l512_id4_0_0_wenable),
    .ram_w16_l512_id4_0_0_enable(ram_w16_l512_id4_0_0_enable),
    .ram_w16_l512_id4_0_1_addr(ram_w16_l512_id4_0_1_addr),
    .ram_w16_l512_id4_0_1_rdata(ram_w16_l512_id4_0_1_rdata),
    .ram_w16_l512_id4_0_1_wdata(ram_w16_l512_id4_0_1_wdata),
    .ram_w16_l512_id4_0_1_wenable(ram_w16_l512_id4_0_1_wenable),
    .ram_w16_l512_id4_0_1_enable(ram_w16_l512_id4_0_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id4_1_0_addr;
  wire [16-1:0] ram_w16_l512_id4_1_0_rdata;
  wire [16-1:0] ram_w16_l512_id4_1_0_wdata;
  wire ram_w16_l512_id4_1_0_wenable;
  wire ram_w16_l512_id4_1_0_enable;
  wire [8-1:0] ram_w16_l512_id4_1_1_addr;
  wire [16-1:0] ram_w16_l512_id4_1_1_rdata;
  wire [16-1:0] ram_w16_l512_id4_1_1_wdata;
  wire ram_w16_l512_id4_1_1_wenable;
  wire ram_w16_l512_id4_1_1_enable;
  assign ram_w16_l512_id4_1_0_wdata = 'hx;
  assign ram_w16_l512_id4_1_0_wenable = 0;

  ram_w16_l512_id4_1
  inst_ram_w16_l512_id4_1
  (
    .CLK(CLK),
    .ram_w16_l512_id4_1_0_addr(ram_w16_l512_id4_1_0_addr),
    .ram_w16_l512_id4_1_0_rdata(ram_w16_l512_id4_1_0_rdata),
    .ram_w16_l512_id4_1_0_wdata(ram_w16_l512_id4_1_0_wdata),
    .ram_w16_l512_id4_1_0_wenable(ram_w16_l512_id4_1_0_wenable),
    .ram_w16_l512_id4_1_0_enable(ram_w16_l512_id4_1_0_enable),
    .ram_w16_l512_id4_1_1_addr(ram_w16_l512_id4_1_1_addr),
    .ram_w16_l512_id4_1_1_rdata(ram_w16_l512_id4_1_1_rdata),
    .ram_w16_l512_id4_1_1_wdata(ram_w16_l512_id4_1_1_wdata),
    .ram_w16_l512_id4_1_1_wenable(ram_w16_l512_id4_1_1_wenable),
    .ram_w16_l512_id4_1_1_enable(ram_w16_l512_id4_1_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id5_0_0_addr;
  wire [16-1:0] ram_w16_l512_id5_0_0_rdata;
  wire [16-1:0] ram_w16_l512_id5_0_0_wdata;
  wire ram_w16_l512_id5_0_0_wenable;
  wire ram_w16_l512_id5_0_0_enable;
  wire [8-1:0] ram_w16_l512_id5_0_1_addr;
  wire [16-1:0] ram_w16_l512_id5_0_1_rdata;
  wire [16-1:0] ram_w16_l512_id5_0_1_wdata;
  wire ram_w16_l512_id5_0_1_wenable;
  wire ram_w16_l512_id5_0_1_enable;
  assign ram_w16_l512_id5_0_0_wdata = 'hx;
  assign ram_w16_l512_id5_0_0_wenable = 0;

  ram_w16_l512_id5_0
  inst_ram_w16_l512_id5_0
  (
    .CLK(CLK),
    .ram_w16_l512_id5_0_0_addr(ram_w16_l512_id5_0_0_addr),
    .ram_w16_l512_id5_0_0_rdata(ram_w16_l512_id5_0_0_rdata),
    .ram_w16_l512_id5_0_0_wdata(ram_w16_l512_id5_0_0_wdata),
    .ram_w16_l512_id5_0_0_wenable(ram_w16_l512_id5_0_0_wenable),
    .ram_w16_l512_id5_0_0_enable(ram_w16_l512_id5_0_0_enable),
    .ram_w16_l512_id5_0_1_addr(ram_w16_l512_id5_0_1_addr),
    .ram_w16_l512_id5_0_1_rdata(ram_w16_l512_id5_0_1_rdata),
    .ram_w16_l512_id5_0_1_wdata(ram_w16_l512_id5_0_1_wdata),
    .ram_w16_l512_id5_0_1_wenable(ram_w16_l512_id5_0_1_wenable),
    .ram_w16_l512_id5_0_1_enable(ram_w16_l512_id5_0_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id5_1_0_addr;
  wire [16-1:0] ram_w16_l512_id5_1_0_rdata;
  wire [16-1:0] ram_w16_l512_id5_1_0_wdata;
  wire ram_w16_l512_id5_1_0_wenable;
  wire ram_w16_l512_id5_1_0_enable;
  wire [8-1:0] ram_w16_l512_id5_1_1_addr;
  wire [16-1:0] ram_w16_l512_id5_1_1_rdata;
  wire [16-1:0] ram_w16_l512_id5_1_1_wdata;
  wire ram_w16_l512_id5_1_1_wenable;
  wire ram_w16_l512_id5_1_1_enable;
  assign ram_w16_l512_id5_1_0_wdata = 'hx;
  assign ram_w16_l512_id5_1_0_wenable = 0;

  ram_w16_l512_id5_1
  inst_ram_w16_l512_id5_1
  (
    .CLK(CLK),
    .ram_w16_l512_id5_1_0_addr(ram_w16_l512_id5_1_0_addr),
    .ram_w16_l512_id5_1_0_rdata(ram_w16_l512_id5_1_0_rdata),
    .ram_w16_l512_id5_1_0_wdata(ram_w16_l512_id5_1_0_wdata),
    .ram_w16_l512_id5_1_0_wenable(ram_w16_l512_id5_1_0_wenable),
    .ram_w16_l512_id5_1_0_enable(ram_w16_l512_id5_1_0_enable),
    .ram_w16_l512_id5_1_1_addr(ram_w16_l512_id5_1_1_addr),
    .ram_w16_l512_id5_1_1_rdata(ram_w16_l512_id5_1_1_rdata),
    .ram_w16_l512_id5_1_1_wdata(ram_w16_l512_id5_1_1_wdata),
    .ram_w16_l512_id5_1_1_wenable(ram_w16_l512_id5_1_1_wenable),
    .ram_w16_l512_id5_1_1_enable(ram_w16_l512_id5_1_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id6_0_0_addr;
  wire [16-1:0] ram_w16_l512_id6_0_0_rdata;
  wire [16-1:0] ram_w16_l512_id6_0_0_wdata;
  wire ram_w16_l512_id6_0_0_wenable;
  wire ram_w16_l512_id6_0_0_enable;
  wire [8-1:0] ram_w16_l512_id6_0_1_addr;
  wire [16-1:0] ram_w16_l512_id6_0_1_rdata;
  wire [16-1:0] ram_w16_l512_id6_0_1_wdata;
  wire ram_w16_l512_id6_0_1_wenable;
  wire ram_w16_l512_id6_0_1_enable;
  assign ram_w16_l512_id6_0_0_wdata = 'hx;
  assign ram_w16_l512_id6_0_0_wenable = 0;

  ram_w16_l512_id6_0
  inst_ram_w16_l512_id6_0
  (
    .CLK(CLK),
    .ram_w16_l512_id6_0_0_addr(ram_w16_l512_id6_0_0_addr),
    .ram_w16_l512_id6_0_0_rdata(ram_w16_l512_id6_0_0_rdata),
    .ram_w16_l512_id6_0_0_wdata(ram_w16_l512_id6_0_0_wdata),
    .ram_w16_l512_id6_0_0_wenable(ram_w16_l512_id6_0_0_wenable),
    .ram_w16_l512_id6_0_0_enable(ram_w16_l512_id6_0_0_enable),
    .ram_w16_l512_id6_0_1_addr(ram_w16_l512_id6_0_1_addr),
    .ram_w16_l512_id6_0_1_rdata(ram_w16_l512_id6_0_1_rdata),
    .ram_w16_l512_id6_0_1_wdata(ram_w16_l512_id6_0_1_wdata),
    .ram_w16_l512_id6_0_1_wenable(ram_w16_l512_id6_0_1_wenable),
    .ram_w16_l512_id6_0_1_enable(ram_w16_l512_id6_0_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id6_1_0_addr;
  wire [16-1:0] ram_w16_l512_id6_1_0_rdata;
  wire [16-1:0] ram_w16_l512_id6_1_0_wdata;
  wire ram_w16_l512_id6_1_0_wenable;
  wire ram_w16_l512_id6_1_0_enable;
  wire [8-1:0] ram_w16_l512_id6_1_1_addr;
  wire [16-1:0] ram_w16_l512_id6_1_1_rdata;
  wire [16-1:0] ram_w16_l512_id6_1_1_wdata;
  wire ram_w16_l512_id6_1_1_wenable;
  wire ram_w16_l512_id6_1_1_enable;
  assign ram_w16_l512_id6_1_0_wdata = 'hx;
  assign ram_w16_l512_id6_1_0_wenable = 0;

  ram_w16_l512_id6_1
  inst_ram_w16_l512_id6_1
  (
    .CLK(CLK),
    .ram_w16_l512_id6_1_0_addr(ram_w16_l512_id6_1_0_addr),
    .ram_w16_l512_id6_1_0_rdata(ram_w16_l512_id6_1_0_rdata),
    .ram_w16_l512_id6_1_0_wdata(ram_w16_l512_id6_1_0_wdata),
    .ram_w16_l512_id6_1_0_wenable(ram_w16_l512_id6_1_0_wenable),
    .ram_w16_l512_id6_1_0_enable(ram_w16_l512_id6_1_0_enable),
    .ram_w16_l512_id6_1_1_addr(ram_w16_l512_id6_1_1_addr),
    .ram_w16_l512_id6_1_1_rdata(ram_w16_l512_id6_1_1_rdata),
    .ram_w16_l512_id6_1_1_wdata(ram_w16_l512_id6_1_1_wdata),
    .ram_w16_l512_id6_1_1_wenable(ram_w16_l512_id6_1_1_wenable),
    .ram_w16_l512_id6_1_1_enable(ram_w16_l512_id6_1_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id7_0_0_addr;
  wire [16-1:0] ram_w16_l512_id7_0_0_rdata;
  wire [16-1:0] ram_w16_l512_id7_0_0_wdata;
  wire ram_w16_l512_id7_0_0_wenable;
  wire ram_w16_l512_id7_0_0_enable;
  wire [8-1:0] ram_w16_l512_id7_0_1_addr;
  wire [16-1:0] ram_w16_l512_id7_0_1_rdata;
  wire [16-1:0] ram_w16_l512_id7_0_1_wdata;
  wire ram_w16_l512_id7_0_1_wenable;
  wire ram_w16_l512_id7_0_1_enable;
  assign ram_w16_l512_id7_0_0_wdata = 'hx;
  assign ram_w16_l512_id7_0_0_wenable = 0;

  ram_w16_l512_id7_0
  inst_ram_w16_l512_id7_0
  (
    .CLK(CLK),
    .ram_w16_l512_id7_0_0_addr(ram_w16_l512_id7_0_0_addr),
    .ram_w16_l512_id7_0_0_rdata(ram_w16_l512_id7_0_0_rdata),
    .ram_w16_l512_id7_0_0_wdata(ram_w16_l512_id7_0_0_wdata),
    .ram_w16_l512_id7_0_0_wenable(ram_w16_l512_id7_0_0_wenable),
    .ram_w16_l512_id7_0_0_enable(ram_w16_l512_id7_0_0_enable),
    .ram_w16_l512_id7_0_1_addr(ram_w16_l512_id7_0_1_addr),
    .ram_w16_l512_id7_0_1_rdata(ram_w16_l512_id7_0_1_rdata),
    .ram_w16_l512_id7_0_1_wdata(ram_w16_l512_id7_0_1_wdata),
    .ram_w16_l512_id7_0_1_wenable(ram_w16_l512_id7_0_1_wenable),
    .ram_w16_l512_id7_0_1_enable(ram_w16_l512_id7_0_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id7_1_0_addr;
  wire [16-1:0] ram_w16_l512_id7_1_0_rdata;
  wire [16-1:0] ram_w16_l512_id7_1_0_wdata;
  wire ram_w16_l512_id7_1_0_wenable;
  wire ram_w16_l512_id7_1_0_enable;
  wire [8-1:0] ram_w16_l512_id7_1_1_addr;
  wire [16-1:0] ram_w16_l512_id7_1_1_rdata;
  wire [16-1:0] ram_w16_l512_id7_1_1_wdata;
  wire ram_w16_l512_id7_1_1_wenable;
  wire ram_w16_l512_id7_1_1_enable;
  assign ram_w16_l512_id7_1_0_wdata = 'hx;
  assign ram_w16_l512_id7_1_0_wenable = 0;

  ram_w16_l512_id7_1
  inst_ram_w16_l512_id7_1
  (
    .CLK(CLK),
    .ram_w16_l512_id7_1_0_addr(ram_w16_l512_id7_1_0_addr),
    .ram_w16_l512_id7_1_0_rdata(ram_w16_l512_id7_1_0_rdata),
    .ram_w16_l512_id7_1_0_wdata(ram_w16_l512_id7_1_0_wdata),
    .ram_w16_l512_id7_1_0_wenable(ram_w16_l512_id7_1_0_wenable),
    .ram_w16_l512_id7_1_0_enable(ram_w16_l512_id7_1_0_enable),
    .ram_w16_l512_id7_1_1_addr(ram_w16_l512_id7_1_1_addr),
    .ram_w16_l512_id7_1_1_rdata(ram_w16_l512_id7_1_1_rdata),
    .ram_w16_l512_id7_1_1_wdata(ram_w16_l512_id7_1_1_wdata),
    .ram_w16_l512_id7_1_1_wenable(ram_w16_l512_id7_1_1_wenable),
    .ram_w16_l512_id7_1_1_enable(ram_w16_l512_id7_1_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id8_0_0_addr;
  wire [16-1:0] ram_w16_l512_id8_0_0_rdata;
  wire [16-1:0] ram_w16_l512_id8_0_0_wdata;
  wire ram_w16_l512_id8_0_0_wenable;
  wire ram_w16_l512_id8_0_0_enable;
  wire [8-1:0] ram_w16_l512_id8_0_1_addr;
  wire [16-1:0] ram_w16_l512_id8_0_1_rdata;
  wire [16-1:0] ram_w16_l512_id8_0_1_wdata;
  wire ram_w16_l512_id8_0_1_wenable;
  wire ram_w16_l512_id8_0_1_enable;
  assign ram_w16_l512_id8_0_0_wdata = 'hx;
  assign ram_w16_l512_id8_0_0_wenable = 0;

  ram_w16_l512_id8_0
  inst_ram_w16_l512_id8_0
  (
    .CLK(CLK),
    .ram_w16_l512_id8_0_0_addr(ram_w16_l512_id8_0_0_addr),
    .ram_w16_l512_id8_0_0_rdata(ram_w16_l512_id8_0_0_rdata),
    .ram_w16_l512_id8_0_0_wdata(ram_w16_l512_id8_0_0_wdata),
    .ram_w16_l512_id8_0_0_wenable(ram_w16_l512_id8_0_0_wenable),
    .ram_w16_l512_id8_0_0_enable(ram_w16_l512_id8_0_0_enable),
    .ram_w16_l512_id8_0_1_addr(ram_w16_l512_id8_0_1_addr),
    .ram_w16_l512_id8_0_1_rdata(ram_w16_l512_id8_0_1_rdata),
    .ram_w16_l512_id8_0_1_wdata(ram_w16_l512_id8_0_1_wdata),
    .ram_w16_l512_id8_0_1_wenable(ram_w16_l512_id8_0_1_wenable),
    .ram_w16_l512_id8_0_1_enable(ram_w16_l512_id8_0_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id8_1_0_addr;
  wire [16-1:0] ram_w16_l512_id8_1_0_rdata;
  wire [16-1:0] ram_w16_l512_id8_1_0_wdata;
  wire ram_w16_l512_id8_1_0_wenable;
  wire ram_w16_l512_id8_1_0_enable;
  wire [8-1:0] ram_w16_l512_id8_1_1_addr;
  wire [16-1:0] ram_w16_l512_id8_1_1_rdata;
  wire [16-1:0] ram_w16_l512_id8_1_1_wdata;
  wire ram_w16_l512_id8_1_1_wenable;
  wire ram_w16_l512_id8_1_1_enable;
  assign ram_w16_l512_id8_1_0_wdata = 'hx;
  assign ram_w16_l512_id8_1_0_wenable = 0;

  ram_w16_l512_id8_1
  inst_ram_w16_l512_id8_1
  (
    .CLK(CLK),
    .ram_w16_l512_id8_1_0_addr(ram_w16_l512_id8_1_0_addr),
    .ram_w16_l512_id8_1_0_rdata(ram_w16_l512_id8_1_0_rdata),
    .ram_w16_l512_id8_1_0_wdata(ram_w16_l512_id8_1_0_wdata),
    .ram_w16_l512_id8_1_0_wenable(ram_w16_l512_id8_1_0_wenable),
    .ram_w16_l512_id8_1_0_enable(ram_w16_l512_id8_1_0_enable),
    .ram_w16_l512_id8_1_1_addr(ram_w16_l512_id8_1_1_addr),
    .ram_w16_l512_id8_1_1_rdata(ram_w16_l512_id8_1_1_rdata),
    .ram_w16_l512_id8_1_1_wdata(ram_w16_l512_id8_1_1_wdata),
    .ram_w16_l512_id8_1_1_wenable(ram_w16_l512_id8_1_1_wenable),
    .ram_w16_l512_id8_1_1_enable(ram_w16_l512_id8_1_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id9_0_0_addr;
  wire [16-1:0] ram_w16_l512_id9_0_0_rdata;
  wire [16-1:0] ram_w16_l512_id9_0_0_wdata;
  wire ram_w16_l512_id9_0_0_wenable;
  wire ram_w16_l512_id9_0_0_enable;
  wire [8-1:0] ram_w16_l512_id9_0_1_addr;
  wire [16-1:0] ram_w16_l512_id9_0_1_rdata;
  wire [16-1:0] ram_w16_l512_id9_0_1_wdata;
  wire ram_w16_l512_id9_0_1_wenable;
  wire ram_w16_l512_id9_0_1_enable;
  assign ram_w16_l512_id9_0_0_wdata = 'hx;
  assign ram_w16_l512_id9_0_0_wenable = 0;

  ram_w16_l512_id9_0
  inst_ram_w16_l512_id9_0
  (
    .CLK(CLK),
    .ram_w16_l512_id9_0_0_addr(ram_w16_l512_id9_0_0_addr),
    .ram_w16_l512_id9_0_0_rdata(ram_w16_l512_id9_0_0_rdata),
    .ram_w16_l512_id9_0_0_wdata(ram_w16_l512_id9_0_0_wdata),
    .ram_w16_l512_id9_0_0_wenable(ram_w16_l512_id9_0_0_wenable),
    .ram_w16_l512_id9_0_0_enable(ram_w16_l512_id9_0_0_enable),
    .ram_w16_l512_id9_0_1_addr(ram_w16_l512_id9_0_1_addr),
    .ram_w16_l512_id9_0_1_rdata(ram_w16_l512_id9_0_1_rdata),
    .ram_w16_l512_id9_0_1_wdata(ram_w16_l512_id9_0_1_wdata),
    .ram_w16_l512_id9_0_1_wenable(ram_w16_l512_id9_0_1_wenable),
    .ram_w16_l512_id9_0_1_enable(ram_w16_l512_id9_0_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id9_1_0_addr;
  wire [16-1:0] ram_w16_l512_id9_1_0_rdata;
  wire [16-1:0] ram_w16_l512_id9_1_0_wdata;
  wire ram_w16_l512_id9_1_0_wenable;
  wire ram_w16_l512_id9_1_0_enable;
  wire [8-1:0] ram_w16_l512_id9_1_1_addr;
  wire [16-1:0] ram_w16_l512_id9_1_1_rdata;
  wire [16-1:0] ram_w16_l512_id9_1_1_wdata;
  wire ram_w16_l512_id9_1_1_wenable;
  wire ram_w16_l512_id9_1_1_enable;
  assign ram_w16_l512_id9_1_0_wdata = 'hx;
  assign ram_w16_l512_id9_1_0_wenable = 0;

  ram_w16_l512_id9_1
  inst_ram_w16_l512_id9_1
  (
    .CLK(CLK),
    .ram_w16_l512_id9_1_0_addr(ram_w16_l512_id9_1_0_addr),
    .ram_w16_l512_id9_1_0_rdata(ram_w16_l512_id9_1_0_rdata),
    .ram_w16_l512_id9_1_0_wdata(ram_w16_l512_id9_1_0_wdata),
    .ram_w16_l512_id9_1_0_wenable(ram_w16_l512_id9_1_0_wenable),
    .ram_w16_l512_id9_1_0_enable(ram_w16_l512_id9_1_0_enable),
    .ram_w16_l512_id9_1_1_addr(ram_w16_l512_id9_1_1_addr),
    .ram_w16_l512_id9_1_1_rdata(ram_w16_l512_id9_1_1_rdata),
    .ram_w16_l512_id9_1_1_wdata(ram_w16_l512_id9_1_1_wdata),
    .ram_w16_l512_id9_1_1_wenable(ram_w16_l512_id9_1_1_wenable),
    .ram_w16_l512_id9_1_1_enable(ram_w16_l512_id9_1_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id10_0_0_addr;
  wire [16-1:0] ram_w16_l512_id10_0_0_rdata;
  wire [16-1:0] ram_w16_l512_id10_0_0_wdata;
  wire ram_w16_l512_id10_0_0_wenable;
  wire ram_w16_l512_id10_0_0_enable;
  wire [8-1:0] ram_w16_l512_id10_0_1_addr;
  wire [16-1:0] ram_w16_l512_id10_0_1_rdata;
  wire [16-1:0] ram_w16_l512_id10_0_1_wdata;
  wire ram_w16_l512_id10_0_1_wenable;
  wire ram_w16_l512_id10_0_1_enable;
  assign ram_w16_l512_id10_0_0_wdata = 'hx;
  assign ram_w16_l512_id10_0_0_wenable = 0;

  ram_w16_l512_id10_0
  inst_ram_w16_l512_id10_0
  (
    .CLK(CLK),
    .ram_w16_l512_id10_0_0_addr(ram_w16_l512_id10_0_0_addr),
    .ram_w16_l512_id10_0_0_rdata(ram_w16_l512_id10_0_0_rdata),
    .ram_w16_l512_id10_0_0_wdata(ram_w16_l512_id10_0_0_wdata),
    .ram_w16_l512_id10_0_0_wenable(ram_w16_l512_id10_0_0_wenable),
    .ram_w16_l512_id10_0_0_enable(ram_w16_l512_id10_0_0_enable),
    .ram_w16_l512_id10_0_1_addr(ram_w16_l512_id10_0_1_addr),
    .ram_w16_l512_id10_0_1_rdata(ram_w16_l512_id10_0_1_rdata),
    .ram_w16_l512_id10_0_1_wdata(ram_w16_l512_id10_0_1_wdata),
    .ram_w16_l512_id10_0_1_wenable(ram_w16_l512_id10_0_1_wenable),
    .ram_w16_l512_id10_0_1_enable(ram_w16_l512_id10_0_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id10_1_0_addr;
  wire [16-1:0] ram_w16_l512_id10_1_0_rdata;
  wire [16-1:0] ram_w16_l512_id10_1_0_wdata;
  wire ram_w16_l512_id10_1_0_wenable;
  wire ram_w16_l512_id10_1_0_enable;
  wire [8-1:0] ram_w16_l512_id10_1_1_addr;
  wire [16-1:0] ram_w16_l512_id10_1_1_rdata;
  wire [16-1:0] ram_w16_l512_id10_1_1_wdata;
  wire ram_w16_l512_id10_1_1_wenable;
  wire ram_w16_l512_id10_1_1_enable;
  assign ram_w16_l512_id10_1_0_wdata = 'hx;
  assign ram_w16_l512_id10_1_0_wenable = 0;

  ram_w16_l512_id10_1
  inst_ram_w16_l512_id10_1
  (
    .CLK(CLK),
    .ram_w16_l512_id10_1_0_addr(ram_w16_l512_id10_1_0_addr),
    .ram_w16_l512_id10_1_0_rdata(ram_w16_l512_id10_1_0_rdata),
    .ram_w16_l512_id10_1_0_wdata(ram_w16_l512_id10_1_0_wdata),
    .ram_w16_l512_id10_1_0_wenable(ram_w16_l512_id10_1_0_wenable),
    .ram_w16_l512_id10_1_0_enable(ram_w16_l512_id10_1_0_enable),
    .ram_w16_l512_id10_1_1_addr(ram_w16_l512_id10_1_1_addr),
    .ram_w16_l512_id10_1_1_rdata(ram_w16_l512_id10_1_1_rdata),
    .ram_w16_l512_id10_1_1_wdata(ram_w16_l512_id10_1_1_wdata),
    .ram_w16_l512_id10_1_1_wenable(ram_w16_l512_id10_1_1_wenable),
    .ram_w16_l512_id10_1_1_enable(ram_w16_l512_id10_1_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id11_0_0_addr;
  wire [16-1:0] ram_w16_l512_id11_0_0_rdata;
  wire [16-1:0] ram_w16_l512_id11_0_0_wdata;
  wire ram_w16_l512_id11_0_0_wenable;
  wire ram_w16_l512_id11_0_0_enable;
  wire [8-1:0] ram_w16_l512_id11_0_1_addr;
  wire [16-1:0] ram_w16_l512_id11_0_1_rdata;
  wire [16-1:0] ram_w16_l512_id11_0_1_wdata;
  wire ram_w16_l512_id11_0_1_wenable;
  wire ram_w16_l512_id11_0_1_enable;
  assign ram_w16_l512_id11_0_0_wdata = 'hx;
  assign ram_w16_l512_id11_0_0_wenable = 0;

  ram_w16_l512_id11_0
  inst_ram_w16_l512_id11_0
  (
    .CLK(CLK),
    .ram_w16_l512_id11_0_0_addr(ram_w16_l512_id11_0_0_addr),
    .ram_w16_l512_id11_0_0_rdata(ram_w16_l512_id11_0_0_rdata),
    .ram_w16_l512_id11_0_0_wdata(ram_w16_l512_id11_0_0_wdata),
    .ram_w16_l512_id11_0_0_wenable(ram_w16_l512_id11_0_0_wenable),
    .ram_w16_l512_id11_0_0_enable(ram_w16_l512_id11_0_0_enable),
    .ram_w16_l512_id11_0_1_addr(ram_w16_l512_id11_0_1_addr),
    .ram_w16_l512_id11_0_1_rdata(ram_w16_l512_id11_0_1_rdata),
    .ram_w16_l512_id11_0_1_wdata(ram_w16_l512_id11_0_1_wdata),
    .ram_w16_l512_id11_0_1_wenable(ram_w16_l512_id11_0_1_wenable),
    .ram_w16_l512_id11_0_1_enable(ram_w16_l512_id11_0_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id11_1_0_addr;
  wire [16-1:0] ram_w16_l512_id11_1_0_rdata;
  wire [16-1:0] ram_w16_l512_id11_1_0_wdata;
  wire ram_w16_l512_id11_1_0_wenable;
  wire ram_w16_l512_id11_1_0_enable;
  wire [8-1:0] ram_w16_l512_id11_1_1_addr;
  wire [16-1:0] ram_w16_l512_id11_1_1_rdata;
  wire [16-1:0] ram_w16_l512_id11_1_1_wdata;
  wire ram_w16_l512_id11_1_1_wenable;
  wire ram_w16_l512_id11_1_1_enable;
  assign ram_w16_l512_id11_1_0_wdata = 'hx;
  assign ram_w16_l512_id11_1_0_wenable = 0;

  ram_w16_l512_id11_1
  inst_ram_w16_l512_id11_1
  (
    .CLK(CLK),
    .ram_w16_l512_id11_1_0_addr(ram_w16_l512_id11_1_0_addr),
    .ram_w16_l512_id11_1_0_rdata(ram_w16_l512_id11_1_0_rdata),
    .ram_w16_l512_id11_1_0_wdata(ram_w16_l512_id11_1_0_wdata),
    .ram_w16_l512_id11_1_0_wenable(ram_w16_l512_id11_1_0_wenable),
    .ram_w16_l512_id11_1_0_enable(ram_w16_l512_id11_1_0_enable),
    .ram_w16_l512_id11_1_1_addr(ram_w16_l512_id11_1_1_addr),
    .ram_w16_l512_id11_1_1_rdata(ram_w16_l512_id11_1_1_rdata),
    .ram_w16_l512_id11_1_1_wdata(ram_w16_l512_id11_1_1_wdata),
    .ram_w16_l512_id11_1_1_wenable(ram_w16_l512_id11_1_1_wenable),
    .ram_w16_l512_id11_1_1_enable(ram_w16_l512_id11_1_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id12_0_0_addr;
  wire [16-1:0] ram_w16_l512_id12_0_0_rdata;
  wire [16-1:0] ram_w16_l512_id12_0_0_wdata;
  wire ram_w16_l512_id12_0_0_wenable;
  wire ram_w16_l512_id12_0_0_enable;
  wire [8-1:0] ram_w16_l512_id12_0_1_addr;
  wire [16-1:0] ram_w16_l512_id12_0_1_rdata;
  wire [16-1:0] ram_w16_l512_id12_0_1_wdata;
  wire ram_w16_l512_id12_0_1_wenable;
  wire ram_w16_l512_id12_0_1_enable;
  assign ram_w16_l512_id12_0_0_wdata = 'hx;
  assign ram_w16_l512_id12_0_0_wenable = 0;

  ram_w16_l512_id12_0
  inst_ram_w16_l512_id12_0
  (
    .CLK(CLK),
    .ram_w16_l512_id12_0_0_addr(ram_w16_l512_id12_0_0_addr),
    .ram_w16_l512_id12_0_0_rdata(ram_w16_l512_id12_0_0_rdata),
    .ram_w16_l512_id12_0_0_wdata(ram_w16_l512_id12_0_0_wdata),
    .ram_w16_l512_id12_0_0_wenable(ram_w16_l512_id12_0_0_wenable),
    .ram_w16_l512_id12_0_0_enable(ram_w16_l512_id12_0_0_enable),
    .ram_w16_l512_id12_0_1_addr(ram_w16_l512_id12_0_1_addr),
    .ram_w16_l512_id12_0_1_rdata(ram_w16_l512_id12_0_1_rdata),
    .ram_w16_l512_id12_0_1_wdata(ram_w16_l512_id12_0_1_wdata),
    .ram_w16_l512_id12_0_1_wenable(ram_w16_l512_id12_0_1_wenable),
    .ram_w16_l512_id12_0_1_enable(ram_w16_l512_id12_0_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id12_1_0_addr;
  wire [16-1:0] ram_w16_l512_id12_1_0_rdata;
  wire [16-1:0] ram_w16_l512_id12_1_0_wdata;
  wire ram_w16_l512_id12_1_0_wenable;
  wire ram_w16_l512_id12_1_0_enable;
  wire [8-1:0] ram_w16_l512_id12_1_1_addr;
  wire [16-1:0] ram_w16_l512_id12_1_1_rdata;
  wire [16-1:0] ram_w16_l512_id12_1_1_wdata;
  wire ram_w16_l512_id12_1_1_wenable;
  wire ram_w16_l512_id12_1_1_enable;
  assign ram_w16_l512_id12_1_0_wdata = 'hx;
  assign ram_w16_l512_id12_1_0_wenable = 0;

  ram_w16_l512_id12_1
  inst_ram_w16_l512_id12_1
  (
    .CLK(CLK),
    .ram_w16_l512_id12_1_0_addr(ram_w16_l512_id12_1_0_addr),
    .ram_w16_l512_id12_1_0_rdata(ram_w16_l512_id12_1_0_rdata),
    .ram_w16_l512_id12_1_0_wdata(ram_w16_l512_id12_1_0_wdata),
    .ram_w16_l512_id12_1_0_wenable(ram_w16_l512_id12_1_0_wenable),
    .ram_w16_l512_id12_1_0_enable(ram_w16_l512_id12_1_0_enable),
    .ram_w16_l512_id12_1_1_addr(ram_w16_l512_id12_1_1_addr),
    .ram_w16_l512_id12_1_1_rdata(ram_w16_l512_id12_1_1_rdata),
    .ram_w16_l512_id12_1_1_wdata(ram_w16_l512_id12_1_1_wdata),
    .ram_w16_l512_id12_1_1_wenable(ram_w16_l512_id12_1_1_wenable),
    .ram_w16_l512_id12_1_1_enable(ram_w16_l512_id12_1_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id13_0_0_addr;
  wire [16-1:0] ram_w16_l512_id13_0_0_rdata;
  wire [16-1:0] ram_w16_l512_id13_0_0_wdata;
  wire ram_w16_l512_id13_0_0_wenable;
  wire ram_w16_l512_id13_0_0_enable;
  wire [8-1:0] ram_w16_l512_id13_0_1_addr;
  wire [16-1:0] ram_w16_l512_id13_0_1_rdata;
  wire [16-1:0] ram_w16_l512_id13_0_1_wdata;
  wire ram_w16_l512_id13_0_1_wenable;
  wire ram_w16_l512_id13_0_1_enable;
  assign ram_w16_l512_id13_0_0_wdata = 'hx;
  assign ram_w16_l512_id13_0_0_wenable = 0;

  ram_w16_l512_id13_0
  inst_ram_w16_l512_id13_0
  (
    .CLK(CLK),
    .ram_w16_l512_id13_0_0_addr(ram_w16_l512_id13_0_0_addr),
    .ram_w16_l512_id13_0_0_rdata(ram_w16_l512_id13_0_0_rdata),
    .ram_w16_l512_id13_0_0_wdata(ram_w16_l512_id13_0_0_wdata),
    .ram_w16_l512_id13_0_0_wenable(ram_w16_l512_id13_0_0_wenable),
    .ram_w16_l512_id13_0_0_enable(ram_w16_l512_id13_0_0_enable),
    .ram_w16_l512_id13_0_1_addr(ram_w16_l512_id13_0_1_addr),
    .ram_w16_l512_id13_0_1_rdata(ram_w16_l512_id13_0_1_rdata),
    .ram_w16_l512_id13_0_1_wdata(ram_w16_l512_id13_0_1_wdata),
    .ram_w16_l512_id13_0_1_wenable(ram_w16_l512_id13_0_1_wenable),
    .ram_w16_l512_id13_0_1_enable(ram_w16_l512_id13_0_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id13_1_0_addr;
  wire [16-1:0] ram_w16_l512_id13_1_0_rdata;
  wire [16-1:0] ram_w16_l512_id13_1_0_wdata;
  wire ram_w16_l512_id13_1_0_wenable;
  wire ram_w16_l512_id13_1_0_enable;
  wire [8-1:0] ram_w16_l512_id13_1_1_addr;
  wire [16-1:0] ram_w16_l512_id13_1_1_rdata;
  wire [16-1:0] ram_w16_l512_id13_1_1_wdata;
  wire ram_w16_l512_id13_1_1_wenable;
  wire ram_w16_l512_id13_1_1_enable;
  assign ram_w16_l512_id13_1_0_wdata = 'hx;
  assign ram_w16_l512_id13_1_0_wenable = 0;

  ram_w16_l512_id13_1
  inst_ram_w16_l512_id13_1
  (
    .CLK(CLK),
    .ram_w16_l512_id13_1_0_addr(ram_w16_l512_id13_1_0_addr),
    .ram_w16_l512_id13_1_0_rdata(ram_w16_l512_id13_1_0_rdata),
    .ram_w16_l512_id13_1_0_wdata(ram_w16_l512_id13_1_0_wdata),
    .ram_w16_l512_id13_1_0_wenable(ram_w16_l512_id13_1_0_wenable),
    .ram_w16_l512_id13_1_0_enable(ram_w16_l512_id13_1_0_enable),
    .ram_w16_l512_id13_1_1_addr(ram_w16_l512_id13_1_1_addr),
    .ram_w16_l512_id13_1_1_rdata(ram_w16_l512_id13_1_1_rdata),
    .ram_w16_l512_id13_1_1_wdata(ram_w16_l512_id13_1_1_wdata),
    .ram_w16_l512_id13_1_1_wenable(ram_w16_l512_id13_1_1_wenable),
    .ram_w16_l512_id13_1_1_enable(ram_w16_l512_id13_1_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id14_0_0_addr;
  wire [16-1:0] ram_w16_l512_id14_0_0_rdata;
  wire [16-1:0] ram_w16_l512_id14_0_0_wdata;
  wire ram_w16_l512_id14_0_0_wenable;
  wire ram_w16_l512_id14_0_0_enable;
  wire [8-1:0] ram_w16_l512_id14_0_1_addr;
  wire [16-1:0] ram_w16_l512_id14_0_1_rdata;
  wire [16-1:0] ram_w16_l512_id14_0_1_wdata;
  wire ram_w16_l512_id14_0_1_wenable;
  wire ram_w16_l512_id14_0_1_enable;
  assign ram_w16_l512_id14_0_0_wdata = 'hx;
  assign ram_w16_l512_id14_0_0_wenable = 0;

  ram_w16_l512_id14_0
  inst_ram_w16_l512_id14_0
  (
    .CLK(CLK),
    .ram_w16_l512_id14_0_0_addr(ram_w16_l512_id14_0_0_addr),
    .ram_w16_l512_id14_0_0_rdata(ram_w16_l512_id14_0_0_rdata),
    .ram_w16_l512_id14_0_0_wdata(ram_w16_l512_id14_0_0_wdata),
    .ram_w16_l512_id14_0_0_wenable(ram_w16_l512_id14_0_0_wenable),
    .ram_w16_l512_id14_0_0_enable(ram_w16_l512_id14_0_0_enable),
    .ram_w16_l512_id14_0_1_addr(ram_w16_l512_id14_0_1_addr),
    .ram_w16_l512_id14_0_1_rdata(ram_w16_l512_id14_0_1_rdata),
    .ram_w16_l512_id14_0_1_wdata(ram_w16_l512_id14_0_1_wdata),
    .ram_w16_l512_id14_0_1_wenable(ram_w16_l512_id14_0_1_wenable),
    .ram_w16_l512_id14_0_1_enable(ram_w16_l512_id14_0_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id14_1_0_addr;
  wire [16-1:0] ram_w16_l512_id14_1_0_rdata;
  wire [16-1:0] ram_w16_l512_id14_1_0_wdata;
  wire ram_w16_l512_id14_1_0_wenable;
  wire ram_w16_l512_id14_1_0_enable;
  wire [8-1:0] ram_w16_l512_id14_1_1_addr;
  wire [16-1:0] ram_w16_l512_id14_1_1_rdata;
  wire [16-1:0] ram_w16_l512_id14_1_1_wdata;
  wire ram_w16_l512_id14_1_1_wenable;
  wire ram_w16_l512_id14_1_1_enable;
  assign ram_w16_l512_id14_1_0_wdata = 'hx;
  assign ram_w16_l512_id14_1_0_wenable = 0;

  ram_w16_l512_id14_1
  inst_ram_w16_l512_id14_1
  (
    .CLK(CLK),
    .ram_w16_l512_id14_1_0_addr(ram_w16_l512_id14_1_0_addr),
    .ram_w16_l512_id14_1_0_rdata(ram_w16_l512_id14_1_0_rdata),
    .ram_w16_l512_id14_1_0_wdata(ram_w16_l512_id14_1_0_wdata),
    .ram_w16_l512_id14_1_0_wenable(ram_w16_l512_id14_1_0_wenable),
    .ram_w16_l512_id14_1_0_enable(ram_w16_l512_id14_1_0_enable),
    .ram_w16_l512_id14_1_1_addr(ram_w16_l512_id14_1_1_addr),
    .ram_w16_l512_id14_1_1_rdata(ram_w16_l512_id14_1_1_rdata),
    .ram_w16_l512_id14_1_1_wdata(ram_w16_l512_id14_1_1_wdata),
    .ram_w16_l512_id14_1_1_wenable(ram_w16_l512_id14_1_1_wenable),
    .ram_w16_l512_id14_1_1_enable(ram_w16_l512_id14_1_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id15_0_0_addr;
  wire [16-1:0] ram_w16_l512_id15_0_0_rdata;
  wire [16-1:0] ram_w16_l512_id15_0_0_wdata;
  wire ram_w16_l512_id15_0_0_wenable;
  wire ram_w16_l512_id15_0_0_enable;
  wire [8-1:0] ram_w16_l512_id15_0_1_addr;
  wire [16-1:0] ram_w16_l512_id15_0_1_rdata;
  wire [16-1:0] ram_w16_l512_id15_0_1_wdata;
  wire ram_w16_l512_id15_0_1_wenable;
  wire ram_w16_l512_id15_0_1_enable;
  assign ram_w16_l512_id15_0_0_wdata = 'hx;
  assign ram_w16_l512_id15_0_0_wenable = 0;

  ram_w16_l512_id15_0
  inst_ram_w16_l512_id15_0
  (
    .CLK(CLK),
    .ram_w16_l512_id15_0_0_addr(ram_w16_l512_id15_0_0_addr),
    .ram_w16_l512_id15_0_0_rdata(ram_w16_l512_id15_0_0_rdata),
    .ram_w16_l512_id15_0_0_wdata(ram_w16_l512_id15_0_0_wdata),
    .ram_w16_l512_id15_0_0_wenable(ram_w16_l512_id15_0_0_wenable),
    .ram_w16_l512_id15_0_0_enable(ram_w16_l512_id15_0_0_enable),
    .ram_w16_l512_id15_0_1_addr(ram_w16_l512_id15_0_1_addr),
    .ram_w16_l512_id15_0_1_rdata(ram_w16_l512_id15_0_1_rdata),
    .ram_w16_l512_id15_0_1_wdata(ram_w16_l512_id15_0_1_wdata),
    .ram_w16_l512_id15_0_1_wenable(ram_w16_l512_id15_0_1_wenable),
    .ram_w16_l512_id15_0_1_enable(ram_w16_l512_id15_0_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id15_1_0_addr;
  wire [16-1:0] ram_w16_l512_id15_1_0_rdata;
  wire [16-1:0] ram_w16_l512_id15_1_0_wdata;
  wire ram_w16_l512_id15_1_0_wenable;
  wire ram_w16_l512_id15_1_0_enable;
  wire [8-1:0] ram_w16_l512_id15_1_1_addr;
  wire [16-1:0] ram_w16_l512_id15_1_1_rdata;
  wire [16-1:0] ram_w16_l512_id15_1_1_wdata;
  wire ram_w16_l512_id15_1_1_wenable;
  wire ram_w16_l512_id15_1_1_enable;
  assign ram_w16_l512_id15_1_0_wdata = 'hx;
  assign ram_w16_l512_id15_1_0_wenable = 0;

  ram_w16_l512_id15_1
  inst_ram_w16_l512_id15_1
  (
    .CLK(CLK),
    .ram_w16_l512_id15_1_0_addr(ram_w16_l512_id15_1_0_addr),
    .ram_w16_l512_id15_1_0_rdata(ram_w16_l512_id15_1_0_rdata),
    .ram_w16_l512_id15_1_0_wdata(ram_w16_l512_id15_1_0_wdata),
    .ram_w16_l512_id15_1_0_wenable(ram_w16_l512_id15_1_0_wenable),
    .ram_w16_l512_id15_1_0_enable(ram_w16_l512_id15_1_0_enable),
    .ram_w16_l512_id15_1_1_addr(ram_w16_l512_id15_1_1_addr),
    .ram_w16_l512_id15_1_1_rdata(ram_w16_l512_id15_1_1_rdata),
    .ram_w16_l512_id15_1_1_wdata(ram_w16_l512_id15_1_1_wdata),
    .ram_w16_l512_id15_1_1_wenable(ram_w16_l512_id15_1_1_wenable),
    .ram_w16_l512_id15_1_1_enable(ram_w16_l512_id15_1_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id16_0_0_addr;
  wire [16-1:0] ram_w16_l512_id16_0_0_rdata;
  wire [16-1:0] ram_w16_l512_id16_0_0_wdata;
  wire ram_w16_l512_id16_0_0_wenable;
  wire ram_w16_l512_id16_0_0_enable;
  wire [8-1:0] ram_w16_l512_id16_0_1_addr;
  wire [16-1:0] ram_w16_l512_id16_0_1_rdata;
  wire [16-1:0] ram_w16_l512_id16_0_1_wdata;
  wire ram_w16_l512_id16_0_1_wenable;
  wire ram_w16_l512_id16_0_1_enable;
  assign ram_w16_l512_id16_0_0_wdata = 'hx;
  assign ram_w16_l512_id16_0_0_wenable = 0;

  ram_w16_l512_id16_0
  inst_ram_w16_l512_id16_0
  (
    .CLK(CLK),
    .ram_w16_l512_id16_0_0_addr(ram_w16_l512_id16_0_0_addr),
    .ram_w16_l512_id16_0_0_rdata(ram_w16_l512_id16_0_0_rdata),
    .ram_w16_l512_id16_0_0_wdata(ram_w16_l512_id16_0_0_wdata),
    .ram_w16_l512_id16_0_0_wenable(ram_w16_l512_id16_0_0_wenable),
    .ram_w16_l512_id16_0_0_enable(ram_w16_l512_id16_0_0_enable),
    .ram_w16_l512_id16_0_1_addr(ram_w16_l512_id16_0_1_addr),
    .ram_w16_l512_id16_0_1_rdata(ram_w16_l512_id16_0_1_rdata),
    .ram_w16_l512_id16_0_1_wdata(ram_w16_l512_id16_0_1_wdata),
    .ram_w16_l512_id16_0_1_wenable(ram_w16_l512_id16_0_1_wenable),
    .ram_w16_l512_id16_0_1_enable(ram_w16_l512_id16_0_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id16_1_0_addr;
  wire [16-1:0] ram_w16_l512_id16_1_0_rdata;
  wire [16-1:0] ram_w16_l512_id16_1_0_wdata;
  wire ram_w16_l512_id16_1_0_wenable;
  wire ram_w16_l512_id16_1_0_enable;
  wire [8-1:0] ram_w16_l512_id16_1_1_addr;
  wire [16-1:0] ram_w16_l512_id16_1_1_rdata;
  wire [16-1:0] ram_w16_l512_id16_1_1_wdata;
  wire ram_w16_l512_id16_1_1_wenable;
  wire ram_w16_l512_id16_1_1_enable;
  assign ram_w16_l512_id16_1_0_wdata = 'hx;
  assign ram_w16_l512_id16_1_0_wenable = 0;

  ram_w16_l512_id16_1
  inst_ram_w16_l512_id16_1
  (
    .CLK(CLK),
    .ram_w16_l512_id16_1_0_addr(ram_w16_l512_id16_1_0_addr),
    .ram_w16_l512_id16_1_0_rdata(ram_w16_l512_id16_1_0_rdata),
    .ram_w16_l512_id16_1_0_wdata(ram_w16_l512_id16_1_0_wdata),
    .ram_w16_l512_id16_1_0_wenable(ram_w16_l512_id16_1_0_wenable),
    .ram_w16_l512_id16_1_0_enable(ram_w16_l512_id16_1_0_enable),
    .ram_w16_l512_id16_1_1_addr(ram_w16_l512_id16_1_1_addr),
    .ram_w16_l512_id16_1_1_rdata(ram_w16_l512_id16_1_1_rdata),
    .ram_w16_l512_id16_1_1_wdata(ram_w16_l512_id16_1_1_wdata),
    .ram_w16_l512_id16_1_1_wenable(ram_w16_l512_id16_1_1_wenable),
    .ram_w16_l512_id16_1_1_enable(ram_w16_l512_id16_1_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id17_0_0_addr;
  wire [16-1:0] ram_w16_l512_id17_0_0_rdata;
  wire [16-1:0] ram_w16_l512_id17_0_0_wdata;
  wire ram_w16_l512_id17_0_0_wenable;
  wire ram_w16_l512_id17_0_0_enable;
  wire [8-1:0] ram_w16_l512_id17_0_1_addr;
  wire [16-1:0] ram_w16_l512_id17_0_1_rdata;
  wire [16-1:0] ram_w16_l512_id17_0_1_wdata;
  wire ram_w16_l512_id17_0_1_wenable;
  wire ram_w16_l512_id17_0_1_enable;
  assign ram_w16_l512_id17_0_0_wdata = 'hx;
  assign ram_w16_l512_id17_0_0_wenable = 0;

  ram_w16_l512_id17_0
  inst_ram_w16_l512_id17_0
  (
    .CLK(CLK),
    .ram_w16_l512_id17_0_0_addr(ram_w16_l512_id17_0_0_addr),
    .ram_w16_l512_id17_0_0_rdata(ram_w16_l512_id17_0_0_rdata),
    .ram_w16_l512_id17_0_0_wdata(ram_w16_l512_id17_0_0_wdata),
    .ram_w16_l512_id17_0_0_wenable(ram_w16_l512_id17_0_0_wenable),
    .ram_w16_l512_id17_0_0_enable(ram_w16_l512_id17_0_0_enable),
    .ram_w16_l512_id17_0_1_addr(ram_w16_l512_id17_0_1_addr),
    .ram_w16_l512_id17_0_1_rdata(ram_w16_l512_id17_0_1_rdata),
    .ram_w16_l512_id17_0_1_wdata(ram_w16_l512_id17_0_1_wdata),
    .ram_w16_l512_id17_0_1_wenable(ram_w16_l512_id17_0_1_wenable),
    .ram_w16_l512_id17_0_1_enable(ram_w16_l512_id17_0_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id17_1_0_addr;
  wire [16-1:0] ram_w16_l512_id17_1_0_rdata;
  wire [16-1:0] ram_w16_l512_id17_1_0_wdata;
  wire ram_w16_l512_id17_1_0_wenable;
  wire ram_w16_l512_id17_1_0_enable;
  wire [8-1:0] ram_w16_l512_id17_1_1_addr;
  wire [16-1:0] ram_w16_l512_id17_1_1_rdata;
  wire [16-1:0] ram_w16_l512_id17_1_1_wdata;
  wire ram_w16_l512_id17_1_1_wenable;
  wire ram_w16_l512_id17_1_1_enable;
  assign ram_w16_l512_id17_1_0_wdata = 'hx;
  assign ram_w16_l512_id17_1_0_wenable = 0;

  ram_w16_l512_id17_1
  inst_ram_w16_l512_id17_1
  (
    .CLK(CLK),
    .ram_w16_l512_id17_1_0_addr(ram_w16_l512_id17_1_0_addr),
    .ram_w16_l512_id17_1_0_rdata(ram_w16_l512_id17_1_0_rdata),
    .ram_w16_l512_id17_1_0_wdata(ram_w16_l512_id17_1_0_wdata),
    .ram_w16_l512_id17_1_0_wenable(ram_w16_l512_id17_1_0_wenable),
    .ram_w16_l512_id17_1_0_enable(ram_w16_l512_id17_1_0_enable),
    .ram_w16_l512_id17_1_1_addr(ram_w16_l512_id17_1_1_addr),
    .ram_w16_l512_id17_1_1_rdata(ram_w16_l512_id17_1_1_rdata),
    .ram_w16_l512_id17_1_1_wdata(ram_w16_l512_id17_1_1_wdata),
    .ram_w16_l512_id17_1_1_wenable(ram_w16_l512_id17_1_1_wenable),
    .ram_w16_l512_id17_1_1_enable(ram_w16_l512_id17_1_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id18_0_0_addr;
  wire [16-1:0] ram_w16_l512_id18_0_0_rdata;
  wire [16-1:0] ram_w16_l512_id18_0_0_wdata;
  wire ram_w16_l512_id18_0_0_wenable;
  wire ram_w16_l512_id18_0_0_enable;
  wire [8-1:0] ram_w16_l512_id18_0_1_addr;
  wire [16-1:0] ram_w16_l512_id18_0_1_rdata;
  wire [16-1:0] ram_w16_l512_id18_0_1_wdata;
  wire ram_w16_l512_id18_0_1_wenable;
  wire ram_w16_l512_id18_0_1_enable;
  assign ram_w16_l512_id18_0_0_wdata = 'hx;
  assign ram_w16_l512_id18_0_0_wenable = 0;

  ram_w16_l512_id18_0
  inst_ram_w16_l512_id18_0
  (
    .CLK(CLK),
    .ram_w16_l512_id18_0_0_addr(ram_w16_l512_id18_0_0_addr),
    .ram_w16_l512_id18_0_0_rdata(ram_w16_l512_id18_0_0_rdata),
    .ram_w16_l512_id18_0_0_wdata(ram_w16_l512_id18_0_0_wdata),
    .ram_w16_l512_id18_0_0_wenable(ram_w16_l512_id18_0_0_wenable),
    .ram_w16_l512_id18_0_0_enable(ram_w16_l512_id18_0_0_enable),
    .ram_w16_l512_id18_0_1_addr(ram_w16_l512_id18_0_1_addr),
    .ram_w16_l512_id18_0_1_rdata(ram_w16_l512_id18_0_1_rdata),
    .ram_w16_l512_id18_0_1_wdata(ram_w16_l512_id18_0_1_wdata),
    .ram_w16_l512_id18_0_1_wenable(ram_w16_l512_id18_0_1_wenable),
    .ram_w16_l512_id18_0_1_enable(ram_w16_l512_id18_0_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id18_1_0_addr;
  wire [16-1:0] ram_w16_l512_id18_1_0_rdata;
  wire [16-1:0] ram_w16_l512_id18_1_0_wdata;
  wire ram_w16_l512_id18_1_0_wenable;
  wire ram_w16_l512_id18_1_0_enable;
  wire [8-1:0] ram_w16_l512_id18_1_1_addr;
  wire [16-1:0] ram_w16_l512_id18_1_1_rdata;
  wire [16-1:0] ram_w16_l512_id18_1_1_wdata;
  wire ram_w16_l512_id18_1_1_wenable;
  wire ram_w16_l512_id18_1_1_enable;
  assign ram_w16_l512_id18_1_0_wdata = 'hx;
  assign ram_w16_l512_id18_1_0_wenable = 0;

  ram_w16_l512_id18_1
  inst_ram_w16_l512_id18_1
  (
    .CLK(CLK),
    .ram_w16_l512_id18_1_0_addr(ram_w16_l512_id18_1_0_addr),
    .ram_w16_l512_id18_1_0_rdata(ram_w16_l512_id18_1_0_rdata),
    .ram_w16_l512_id18_1_0_wdata(ram_w16_l512_id18_1_0_wdata),
    .ram_w16_l512_id18_1_0_wenable(ram_w16_l512_id18_1_0_wenable),
    .ram_w16_l512_id18_1_0_enable(ram_w16_l512_id18_1_0_enable),
    .ram_w16_l512_id18_1_1_addr(ram_w16_l512_id18_1_1_addr),
    .ram_w16_l512_id18_1_1_rdata(ram_w16_l512_id18_1_1_rdata),
    .ram_w16_l512_id18_1_1_wdata(ram_w16_l512_id18_1_1_wdata),
    .ram_w16_l512_id18_1_1_wenable(ram_w16_l512_id18_1_1_wenable),
    .ram_w16_l512_id18_1_1_enable(ram_w16_l512_id18_1_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id19_0_0_addr;
  wire [16-1:0] ram_w16_l512_id19_0_0_rdata;
  wire [16-1:0] ram_w16_l512_id19_0_0_wdata;
  wire ram_w16_l512_id19_0_0_wenable;
  wire ram_w16_l512_id19_0_0_enable;
  wire [8-1:0] ram_w16_l512_id19_0_1_addr;
  wire [16-1:0] ram_w16_l512_id19_0_1_rdata;
  wire [16-1:0] ram_w16_l512_id19_0_1_wdata;
  wire ram_w16_l512_id19_0_1_wenable;
  wire ram_w16_l512_id19_0_1_enable;
  assign ram_w16_l512_id19_0_0_wdata = 'hx;
  assign ram_w16_l512_id19_0_0_wenable = 0;

  ram_w16_l512_id19_0
  inst_ram_w16_l512_id19_0
  (
    .CLK(CLK),
    .ram_w16_l512_id19_0_0_addr(ram_w16_l512_id19_0_0_addr),
    .ram_w16_l512_id19_0_0_rdata(ram_w16_l512_id19_0_0_rdata),
    .ram_w16_l512_id19_0_0_wdata(ram_w16_l512_id19_0_0_wdata),
    .ram_w16_l512_id19_0_0_wenable(ram_w16_l512_id19_0_0_wenable),
    .ram_w16_l512_id19_0_0_enable(ram_w16_l512_id19_0_0_enable),
    .ram_w16_l512_id19_0_1_addr(ram_w16_l512_id19_0_1_addr),
    .ram_w16_l512_id19_0_1_rdata(ram_w16_l512_id19_0_1_rdata),
    .ram_w16_l512_id19_0_1_wdata(ram_w16_l512_id19_0_1_wdata),
    .ram_w16_l512_id19_0_1_wenable(ram_w16_l512_id19_0_1_wenable),
    .ram_w16_l512_id19_0_1_enable(ram_w16_l512_id19_0_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id19_1_0_addr;
  wire [16-1:0] ram_w16_l512_id19_1_0_rdata;
  wire [16-1:0] ram_w16_l512_id19_1_0_wdata;
  wire ram_w16_l512_id19_1_0_wenable;
  wire ram_w16_l512_id19_1_0_enable;
  wire [8-1:0] ram_w16_l512_id19_1_1_addr;
  wire [16-1:0] ram_w16_l512_id19_1_1_rdata;
  wire [16-1:0] ram_w16_l512_id19_1_1_wdata;
  wire ram_w16_l512_id19_1_1_wenable;
  wire ram_w16_l512_id19_1_1_enable;
  assign ram_w16_l512_id19_1_0_wdata = 'hx;
  assign ram_w16_l512_id19_1_0_wenable = 0;

  ram_w16_l512_id19_1
  inst_ram_w16_l512_id19_1
  (
    .CLK(CLK),
    .ram_w16_l512_id19_1_0_addr(ram_w16_l512_id19_1_0_addr),
    .ram_w16_l512_id19_1_0_rdata(ram_w16_l512_id19_1_0_rdata),
    .ram_w16_l512_id19_1_0_wdata(ram_w16_l512_id19_1_0_wdata),
    .ram_w16_l512_id19_1_0_wenable(ram_w16_l512_id19_1_0_wenable),
    .ram_w16_l512_id19_1_0_enable(ram_w16_l512_id19_1_0_enable),
    .ram_w16_l512_id19_1_1_addr(ram_w16_l512_id19_1_1_addr),
    .ram_w16_l512_id19_1_1_rdata(ram_w16_l512_id19_1_1_rdata),
    .ram_w16_l512_id19_1_1_wdata(ram_w16_l512_id19_1_1_wdata),
    .ram_w16_l512_id19_1_1_wenable(ram_w16_l512_id19_1_1_wenable),
    .ram_w16_l512_id19_1_1_enable(ram_w16_l512_id19_1_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id20_0_0_addr;
  wire [16-1:0] ram_w16_l512_id20_0_0_rdata;
  wire [16-1:0] ram_w16_l512_id20_0_0_wdata;
  wire ram_w16_l512_id20_0_0_wenable;
  wire ram_w16_l512_id20_0_0_enable;
  wire [8-1:0] ram_w16_l512_id20_0_1_addr;
  wire [16-1:0] ram_w16_l512_id20_0_1_rdata;
  wire [16-1:0] ram_w16_l512_id20_0_1_wdata;
  wire ram_w16_l512_id20_0_1_wenable;
  wire ram_w16_l512_id20_0_1_enable;
  assign ram_w16_l512_id20_0_1_wdata = 'hx;
  assign ram_w16_l512_id20_0_1_wenable = 0;

  ram_w16_l512_id20_0
  inst_ram_w16_l512_id20_0
  (
    .CLK(CLK),
    .ram_w16_l512_id20_0_0_addr(ram_w16_l512_id20_0_0_addr),
    .ram_w16_l512_id20_0_0_rdata(ram_w16_l512_id20_0_0_rdata),
    .ram_w16_l512_id20_0_0_wdata(ram_w16_l512_id20_0_0_wdata),
    .ram_w16_l512_id20_0_0_wenable(ram_w16_l512_id20_0_0_wenable),
    .ram_w16_l512_id20_0_0_enable(ram_w16_l512_id20_0_0_enable),
    .ram_w16_l512_id20_0_1_addr(ram_w16_l512_id20_0_1_addr),
    .ram_w16_l512_id20_0_1_rdata(ram_w16_l512_id20_0_1_rdata),
    .ram_w16_l512_id20_0_1_wdata(ram_w16_l512_id20_0_1_wdata),
    .ram_w16_l512_id20_0_1_wenable(ram_w16_l512_id20_0_1_wenable),
    .ram_w16_l512_id20_0_1_enable(ram_w16_l512_id20_0_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id20_1_0_addr;
  wire [16-1:0] ram_w16_l512_id20_1_0_rdata;
  wire [16-1:0] ram_w16_l512_id20_1_0_wdata;
  wire ram_w16_l512_id20_1_0_wenable;
  wire ram_w16_l512_id20_1_0_enable;
  wire [8-1:0] ram_w16_l512_id20_1_1_addr;
  wire [16-1:0] ram_w16_l512_id20_1_1_rdata;
  wire [16-1:0] ram_w16_l512_id20_1_1_wdata;
  wire ram_w16_l512_id20_1_1_wenable;
  wire ram_w16_l512_id20_1_1_enable;
  assign ram_w16_l512_id20_1_1_wdata = 'hx;
  assign ram_w16_l512_id20_1_1_wenable = 0;

  ram_w16_l512_id20_1
  inst_ram_w16_l512_id20_1
  (
    .CLK(CLK),
    .ram_w16_l512_id20_1_0_addr(ram_w16_l512_id20_1_0_addr),
    .ram_w16_l512_id20_1_0_rdata(ram_w16_l512_id20_1_0_rdata),
    .ram_w16_l512_id20_1_0_wdata(ram_w16_l512_id20_1_0_wdata),
    .ram_w16_l512_id20_1_0_wenable(ram_w16_l512_id20_1_0_wenable),
    .ram_w16_l512_id20_1_0_enable(ram_w16_l512_id20_1_0_enable),
    .ram_w16_l512_id20_1_1_addr(ram_w16_l512_id20_1_1_addr),
    .ram_w16_l512_id20_1_1_rdata(ram_w16_l512_id20_1_1_rdata),
    .ram_w16_l512_id20_1_1_wdata(ram_w16_l512_id20_1_1_wdata),
    .ram_w16_l512_id20_1_1_wenable(ram_w16_l512_id20_1_1_wenable),
    .ram_w16_l512_id20_1_1_enable(ram_w16_l512_id20_1_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id21_0_0_addr;
  wire [16-1:0] ram_w16_l512_id21_0_0_rdata;
  wire [16-1:0] ram_w16_l512_id21_0_0_wdata;
  wire ram_w16_l512_id21_0_0_wenable;
  wire ram_w16_l512_id21_0_0_enable;
  wire [8-1:0] ram_w16_l512_id21_0_1_addr;
  wire [16-1:0] ram_w16_l512_id21_0_1_rdata;
  wire [16-1:0] ram_w16_l512_id21_0_1_wdata;
  wire ram_w16_l512_id21_0_1_wenable;
  wire ram_w16_l512_id21_0_1_enable;
  assign ram_w16_l512_id21_0_0_addr = 'hx;
  assign ram_w16_l512_id21_0_0_wdata = 'hx;
  assign ram_w16_l512_id21_0_0_wenable = 0;
  assign ram_w16_l512_id21_0_0_enable = 0;
  assign ram_w16_l512_id21_0_1_addr = 'hx;
  assign ram_w16_l512_id21_0_1_wdata = 'hx;
  assign ram_w16_l512_id21_0_1_wenable = 0;
  assign ram_w16_l512_id21_0_1_enable = 0;

  ram_w16_l512_id21_0
  inst_ram_w16_l512_id21_0
  (
    .CLK(CLK),
    .ram_w16_l512_id21_0_0_addr(ram_w16_l512_id21_0_0_addr),
    .ram_w16_l512_id21_0_0_rdata(ram_w16_l512_id21_0_0_rdata),
    .ram_w16_l512_id21_0_0_wdata(ram_w16_l512_id21_0_0_wdata),
    .ram_w16_l512_id21_0_0_wenable(ram_w16_l512_id21_0_0_wenable),
    .ram_w16_l512_id21_0_0_enable(ram_w16_l512_id21_0_0_enable),
    .ram_w16_l512_id21_0_1_addr(ram_w16_l512_id21_0_1_addr),
    .ram_w16_l512_id21_0_1_rdata(ram_w16_l512_id21_0_1_rdata),
    .ram_w16_l512_id21_0_1_wdata(ram_w16_l512_id21_0_1_wdata),
    .ram_w16_l512_id21_0_1_wenable(ram_w16_l512_id21_0_1_wenable),
    .ram_w16_l512_id21_0_1_enable(ram_w16_l512_id21_0_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id21_1_0_addr;
  wire [16-1:0] ram_w16_l512_id21_1_0_rdata;
  wire [16-1:0] ram_w16_l512_id21_1_0_wdata;
  wire ram_w16_l512_id21_1_0_wenable;
  wire ram_w16_l512_id21_1_0_enable;
  wire [8-1:0] ram_w16_l512_id21_1_1_addr;
  wire [16-1:0] ram_w16_l512_id21_1_1_rdata;
  wire [16-1:0] ram_w16_l512_id21_1_1_wdata;
  wire ram_w16_l512_id21_1_1_wenable;
  wire ram_w16_l512_id21_1_1_enable;
  assign ram_w16_l512_id21_1_0_addr = 'hx;
  assign ram_w16_l512_id21_1_0_wdata = 'hx;
  assign ram_w16_l512_id21_1_0_wenable = 0;
  assign ram_w16_l512_id21_1_0_enable = 0;
  assign ram_w16_l512_id21_1_1_addr = 'hx;
  assign ram_w16_l512_id21_1_1_wdata = 'hx;
  assign ram_w16_l512_id21_1_1_wenable = 0;
  assign ram_w16_l512_id21_1_1_enable = 0;

  ram_w16_l512_id21_1
  inst_ram_w16_l512_id21_1
  (
    .CLK(CLK),
    .ram_w16_l512_id21_1_0_addr(ram_w16_l512_id21_1_0_addr),
    .ram_w16_l512_id21_1_0_rdata(ram_w16_l512_id21_1_0_rdata),
    .ram_w16_l512_id21_1_0_wdata(ram_w16_l512_id21_1_0_wdata),
    .ram_w16_l512_id21_1_0_wenable(ram_w16_l512_id21_1_0_wenable),
    .ram_w16_l512_id21_1_0_enable(ram_w16_l512_id21_1_0_enable),
    .ram_w16_l512_id21_1_1_addr(ram_w16_l512_id21_1_1_addr),
    .ram_w16_l512_id21_1_1_rdata(ram_w16_l512_id21_1_1_rdata),
    .ram_w16_l512_id21_1_1_wdata(ram_w16_l512_id21_1_1_wdata),
    .ram_w16_l512_id21_1_1_wenable(ram_w16_l512_id21_1_1_wenable),
    .ram_w16_l512_id21_1_1_enable(ram_w16_l512_id21_1_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id22_0_0_addr;
  wire [16-1:0] ram_w16_l512_id22_0_0_rdata;
  wire [16-1:0] ram_w16_l512_id22_0_0_wdata;
  wire ram_w16_l512_id22_0_0_wenable;
  wire ram_w16_l512_id22_0_0_enable;
  wire [8-1:0] ram_w16_l512_id22_0_1_addr;
  wire [16-1:0] ram_w16_l512_id22_0_1_rdata;
  wire [16-1:0] ram_w16_l512_id22_0_1_wdata;
  wire ram_w16_l512_id22_0_1_wenable;
  wire ram_w16_l512_id22_0_1_enable;
  assign ram_w16_l512_id22_0_0_addr = 'hx;
  assign ram_w16_l512_id22_0_0_wdata = 'hx;
  assign ram_w16_l512_id22_0_0_wenable = 0;
  assign ram_w16_l512_id22_0_0_enable = 0;
  assign ram_w16_l512_id22_0_1_addr = 'hx;
  assign ram_w16_l512_id22_0_1_wdata = 'hx;
  assign ram_w16_l512_id22_0_1_wenable = 0;
  assign ram_w16_l512_id22_0_1_enable = 0;

  ram_w16_l512_id22_0
  inst_ram_w16_l512_id22_0
  (
    .CLK(CLK),
    .ram_w16_l512_id22_0_0_addr(ram_w16_l512_id22_0_0_addr),
    .ram_w16_l512_id22_0_0_rdata(ram_w16_l512_id22_0_0_rdata),
    .ram_w16_l512_id22_0_0_wdata(ram_w16_l512_id22_0_0_wdata),
    .ram_w16_l512_id22_0_0_wenable(ram_w16_l512_id22_0_0_wenable),
    .ram_w16_l512_id22_0_0_enable(ram_w16_l512_id22_0_0_enable),
    .ram_w16_l512_id22_0_1_addr(ram_w16_l512_id22_0_1_addr),
    .ram_w16_l512_id22_0_1_rdata(ram_w16_l512_id22_0_1_rdata),
    .ram_w16_l512_id22_0_1_wdata(ram_w16_l512_id22_0_1_wdata),
    .ram_w16_l512_id22_0_1_wenable(ram_w16_l512_id22_0_1_wenable),
    .ram_w16_l512_id22_0_1_enable(ram_w16_l512_id22_0_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id22_1_0_addr;
  wire [16-1:0] ram_w16_l512_id22_1_0_rdata;
  wire [16-1:0] ram_w16_l512_id22_1_0_wdata;
  wire ram_w16_l512_id22_1_0_wenable;
  wire ram_w16_l512_id22_1_0_enable;
  wire [8-1:0] ram_w16_l512_id22_1_1_addr;
  wire [16-1:0] ram_w16_l512_id22_1_1_rdata;
  wire [16-1:0] ram_w16_l512_id22_1_1_wdata;
  wire ram_w16_l512_id22_1_1_wenable;
  wire ram_w16_l512_id22_1_1_enable;
  assign ram_w16_l512_id22_1_0_addr = 'hx;
  assign ram_w16_l512_id22_1_0_wdata = 'hx;
  assign ram_w16_l512_id22_1_0_wenable = 0;
  assign ram_w16_l512_id22_1_0_enable = 0;
  assign ram_w16_l512_id22_1_1_addr = 'hx;
  assign ram_w16_l512_id22_1_1_wdata = 'hx;
  assign ram_w16_l512_id22_1_1_wenable = 0;
  assign ram_w16_l512_id22_1_1_enable = 0;

  ram_w16_l512_id22_1
  inst_ram_w16_l512_id22_1
  (
    .CLK(CLK),
    .ram_w16_l512_id22_1_0_addr(ram_w16_l512_id22_1_0_addr),
    .ram_w16_l512_id22_1_0_rdata(ram_w16_l512_id22_1_0_rdata),
    .ram_w16_l512_id22_1_0_wdata(ram_w16_l512_id22_1_0_wdata),
    .ram_w16_l512_id22_1_0_wenable(ram_w16_l512_id22_1_0_wenable),
    .ram_w16_l512_id22_1_0_enable(ram_w16_l512_id22_1_0_enable),
    .ram_w16_l512_id22_1_1_addr(ram_w16_l512_id22_1_1_addr),
    .ram_w16_l512_id22_1_1_rdata(ram_w16_l512_id22_1_1_rdata),
    .ram_w16_l512_id22_1_1_wdata(ram_w16_l512_id22_1_1_wdata),
    .ram_w16_l512_id22_1_1_wenable(ram_w16_l512_id22_1_1_wenable),
    .ram_w16_l512_id22_1_1_enable(ram_w16_l512_id22_1_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id23_0_0_addr;
  wire [16-1:0] ram_w16_l512_id23_0_0_rdata;
  wire [16-1:0] ram_w16_l512_id23_0_0_wdata;
  wire ram_w16_l512_id23_0_0_wenable;
  wire ram_w16_l512_id23_0_0_enable;
  wire [8-1:0] ram_w16_l512_id23_0_1_addr;
  wire [16-1:0] ram_w16_l512_id23_0_1_rdata;
  wire [16-1:0] ram_w16_l512_id23_0_1_wdata;
  wire ram_w16_l512_id23_0_1_wenable;
  wire ram_w16_l512_id23_0_1_enable;
  assign ram_w16_l512_id23_0_0_addr = 'hx;
  assign ram_w16_l512_id23_0_0_wdata = 'hx;
  assign ram_w16_l512_id23_0_0_wenable = 0;
  assign ram_w16_l512_id23_0_0_enable = 0;
  assign ram_w16_l512_id23_0_1_addr = 'hx;
  assign ram_w16_l512_id23_0_1_wdata = 'hx;
  assign ram_w16_l512_id23_0_1_wenable = 0;
  assign ram_w16_l512_id23_0_1_enable = 0;

  ram_w16_l512_id23_0
  inst_ram_w16_l512_id23_0
  (
    .CLK(CLK),
    .ram_w16_l512_id23_0_0_addr(ram_w16_l512_id23_0_0_addr),
    .ram_w16_l512_id23_0_0_rdata(ram_w16_l512_id23_0_0_rdata),
    .ram_w16_l512_id23_0_0_wdata(ram_w16_l512_id23_0_0_wdata),
    .ram_w16_l512_id23_0_0_wenable(ram_w16_l512_id23_0_0_wenable),
    .ram_w16_l512_id23_0_0_enable(ram_w16_l512_id23_0_0_enable),
    .ram_w16_l512_id23_0_1_addr(ram_w16_l512_id23_0_1_addr),
    .ram_w16_l512_id23_0_1_rdata(ram_w16_l512_id23_0_1_rdata),
    .ram_w16_l512_id23_0_1_wdata(ram_w16_l512_id23_0_1_wdata),
    .ram_w16_l512_id23_0_1_wenable(ram_w16_l512_id23_0_1_wenable),
    .ram_w16_l512_id23_0_1_enable(ram_w16_l512_id23_0_1_enable)
  );

  wire [8-1:0] ram_w16_l512_id23_1_0_addr;
  wire [16-1:0] ram_w16_l512_id23_1_0_rdata;
  wire [16-1:0] ram_w16_l512_id23_1_0_wdata;
  wire ram_w16_l512_id23_1_0_wenable;
  wire ram_w16_l512_id23_1_0_enable;
  wire [8-1:0] ram_w16_l512_id23_1_1_addr;
  wire [16-1:0] ram_w16_l512_id23_1_1_rdata;
  wire [16-1:0] ram_w16_l512_id23_1_1_wdata;
  wire ram_w16_l512_id23_1_1_wenable;
  wire ram_w16_l512_id23_1_1_enable;
  assign ram_w16_l512_id23_1_0_addr = 'hx;
  assign ram_w16_l512_id23_1_0_wdata = 'hx;
  assign ram_w16_l512_id23_1_0_wenable = 0;
  assign ram_w16_l512_id23_1_0_enable = 0;
  assign ram_w16_l512_id23_1_1_addr = 'hx;
  assign ram_w16_l512_id23_1_1_wdata = 'hx;
  assign ram_w16_l512_id23_1_1_wenable = 0;
  assign ram_w16_l512_id23_1_1_enable = 0;

  ram_w16_l512_id23_1
  inst_ram_w16_l512_id23_1
  (
    .CLK(CLK),
    .ram_w16_l512_id23_1_0_addr(ram_w16_l512_id23_1_0_addr),
    .ram_w16_l512_id23_1_0_rdata(ram_w16_l512_id23_1_0_rdata),
    .ram_w16_l512_id23_1_0_wdata(ram_w16_l512_id23_1_0_wdata),
    .ram_w16_l512_id23_1_0_wenable(ram_w16_l512_id23_1_0_wenable),
    .ram_w16_l512_id23_1_0_enable(ram_w16_l512_id23_1_0_enable),
    .ram_w16_l512_id23_1_1_addr(ram_w16_l512_id23_1_1_addr),
    .ram_w16_l512_id23_1_1_rdata(ram_w16_l512_id23_1_1_rdata),
    .ram_w16_l512_id23_1_1_wdata(ram_w16_l512_id23_1_1_wdata),
    .ram_w16_l512_id23_1_1_wenable(ram_w16_l512_id23_1_1_wenable),
    .ram_w16_l512_id23_1_1_enable(ram_w16_l512_id23_1_1_enable)
  );

  wire [5-1:0] cparam_conv2d_4_act_num_col;
  wire [5-1:0] cparam_conv2d_4_act_num_row;
  wire [6-1:0] cparam_conv2d_4_filter_num_och;
  wire [1-1:0] cparam_conv2d_4_bias_scala;
  wire [6-1:0] cparam_conv2d_4_bias_num;
  wire [1-1:0] cparam_conv2d_4_scale_scala;
  wire [6-1:0] cparam_conv2d_4_scale_num;
  wire [1-1:0] cparam_conv2d_4_vshamt_mul_scala;
  wire [1-1:0] cparam_conv2d_4_vshamt_mul_num;
  wire [1-1:0] cparam_conv2d_4_vshamt_sum_scala;
  wire [1-1:0] cparam_conv2d_4_vshamt_sum_num;
  wire [1-1:0] cparam_conv2d_4_vshamt_out_scala;
  wire [1-1:0] cparam_conv2d_4_vshamt_out_num;
  wire [1-1:0] cparam_conv2d_4_cshamt_mul_value;
  wire [1-1:0] cparam_conv2d_4_cshamt_sum_value;
  wire [5-1:0] cparam_conv2d_4_cshamt_out_value;
  wire [1-1:0] cparam_conv2d_4_act_func_index;
  wire [5-1:0] cparam_conv2d_4_out_num_col;
  wire [5-1:0] cparam_conv2d_4_out_num_row;
  wire [1-1:0] cparam_conv2d_4_pad_col_left;
  wire [1-1:0] cparam_conv2d_4_pad_row_top;
  wire [5-1:0] cparam_conv2d_4_max_col_count;
  wire [5-1:0] cparam_conv2d_4_max_row_count;
  wire [1-1:0] cparam_conv2d_4_max_bat_count;
  wire [5-1:0] cparam_conv2d_4_max_och_count;
  wire [4-1:0] cparam_conv2d_4_och_count_step;
  wire [1-1:0] cparam_conv2d_4_dma_flag_conds_0;
  wire [1-1:0] cparam_conv2d_4_dma_flag_conds_1;
  wire [1-1:0] cparam_conv2d_4_dma_flag_conds_2;
  wire signed [32-1:0] cparam_conv2d_4_act_offset_values_0;
  wire signed [32-1:0] cparam_conv2d_4_act_offset_values_1;
  wire signed [32-1:0] cparam_conv2d_4_act_offset_values_2;
  wire [7-1:0] cparam_conv2d_4_act_row_step;
  wire [12-1:0] cparam_conv2d_4_act_bat_step;
  wire [6-1:0] cparam_conv2d_4_act_read_size;
  wire [2-1:0] cparam_conv2d_4_act_read_block;
  wire [5-1:0] cparam_conv2d_4_act_read_step;
  wire [9-1:0] cparam_conv2d_4_filter_base_step;
  wire [8-1:0] cparam_conv2d_4_filter_read_size;
  wire [2-1:0] cparam_conv2d_4_filter_read_block;
  wire [5-1:0] cparam_conv2d_4_filter_read_step;
  wire [1-1:0] cparam_conv2d_4_out_offset_values_0;
  wire [7-1:0] cparam_conv2d_4_out_col_step;
  wire [11-1:0] cparam_conv2d_4_out_row_step;
  wire [16-1:0] cparam_conv2d_4_out_bat_step;
  wire [5-1:0] cparam_conv2d_4_out_och_step;
  wire [4-1:0] cparam_conv2d_4_out_write_size;
  wire [4-1:0] cparam_conv2d_4_out_write_size_res;
  wire [1-1:0] cparam_conv2d_4_out_write_block;
  wire [1-1:0] cparam_conv2d_4_keep_filter;
  wire [1-1:0] cparam_conv2d_4_keep_input;
  wire [1-1:0] cparam_conv2d_4_data_stationary;
  wire [4-1:0] cparam_conv2d_4_stream_num_ops;
  wire [4-1:0] cparam_conv2d_4_stream_num_ops_res;
  wire [4-1:0] cparam_conv2d_4_stream_num_ops_par;
  wire [4-1:0] cparam_conv2d_4_stream_num_ops_res_par;
  wire [1-1:0] cparam_conv2d_4_stream_reduce_size;
  wire [2-1:0] cparam_conv2d_4_stream_aligned_reduce_size;
  wire [1-1:0] cparam_conv2d_4_stream_omit_mask;
  wire [2-1:0] cparam_conv2d_4_col_select_initval;
  wire [1-1:0] cparam_conv2d_4_stride_col_par_col;
  wire [1-1:0] cparam_conv2d_4_stride_row_par_row;
  wire [1-1:0] cparam_conv2d_4_stride_col_mod_filter_num;
  wire [2-1:0] cparam_conv2d_4_filter_num_col_minus_stride_col_mod;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_0;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_1;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_2;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_3;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_4;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_5;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_6;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_7;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_8;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_9;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_10;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_11;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_12;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_13;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_14;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_15;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_16;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_17;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_18;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_19;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_20;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_21;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_22;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_23;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_24;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_25;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_conds_26;
  wire [1-1:0] cparam_conv2d_4_inc_act_laddr_small;
  wire [2-1:0] cparam_conv2d_4_inc_act_laddr_large;
  wire [6-1:0] cparam_conv2d_4_inc_out_laddr_col;
  wire [1-1:0] cparam_conv2d_4_stream_act_local_small_offset;
  wire signed [3-1:0] cparam_conv2d_4_stream_act_local_large_offset;
  wire [1-1:0] cparam_conv2d_4_stream_act_local_small_flags_0;
  wire [1-1:0] cparam_conv2d_4_stream_act_local_small_flags_1;
  wire [1-1:0] cparam_conv2d_4_stream_act_local_small_flags_2;
  wire [1-1:0] cparam_conv2d_4_stream_act_local_large_flags_0;
  wire [1-1:0] cparam_conv2d_4_stream_act_local_large_flags_1;
  wire [1-1:0] cparam_conv2d_4_stream_act_local_large_flags_2;
  wire [1-1:0] cparam_conv2d_4_inc_sync_out;
  wire [1-1:0] cparam_conv2d_4_inc_sync_out_res;
  assign cparam_conv2d_4_act_num_col = 28;
  assign cparam_conv2d_4_act_num_row = 28;
  assign cparam_conv2d_4_filter_num_och = 32;
  assign cparam_conv2d_4_bias_scala = 0;
  assign cparam_conv2d_4_bias_num = 32;
  assign cparam_conv2d_4_scale_scala = 0;
  assign cparam_conv2d_4_scale_num = 32;
  assign cparam_conv2d_4_vshamt_mul_scala = 0;
  assign cparam_conv2d_4_vshamt_mul_num = 0;
  assign cparam_conv2d_4_vshamt_sum_scala = 0;
  assign cparam_conv2d_4_vshamt_sum_num = 0;
  assign cparam_conv2d_4_vshamt_out_scala = 0;
  assign cparam_conv2d_4_vshamt_out_num = 0;
  assign cparam_conv2d_4_cshamt_mul_value = 0;
  assign cparam_conv2d_4_cshamt_sum_value = 0;
  assign cparam_conv2d_4_cshamt_out_value = 30;
  assign cparam_conv2d_4_act_func_index = 0;
  assign cparam_conv2d_4_out_num_col = 28;
  assign cparam_conv2d_4_out_num_row = 28;
  assign cparam_conv2d_4_pad_col_left = 1;
  assign cparam_conv2d_4_pad_row_top = 1;
  assign cparam_conv2d_4_max_col_count = 27;
  assign cparam_conv2d_4_max_row_count = 27;
  assign cparam_conv2d_4_max_bat_count = 0;
  assign cparam_conv2d_4_max_och_count = 24;
  assign cparam_conv2d_4_och_count_step = 8;
  assign cparam_conv2d_4_dma_flag_conds_0 = 1;
  assign cparam_conv2d_4_dma_flag_conds_1 = 0;
  assign cparam_conv2d_4_dma_flag_conds_2 = 0;
  assign cparam_conv2d_4_act_offset_values_0 = -112;
  assign cparam_conv2d_4_act_offset_values_1 = 0;
  assign cparam_conv2d_4_act_offset_values_2 = 112;
  assign cparam_conv2d_4_act_row_step = 112;
  assign cparam_conv2d_4_act_bat_step = 3136;
  assign cparam_conv2d_4_act_read_size = 56;
  assign cparam_conv2d_4_act_read_block = 2;
  assign cparam_conv2d_4_act_read_step = 20;
  assign cparam_conv2d_4_filter_base_step = 288;
  assign cparam_conv2d_4_filter_read_size = 144;
  assign cparam_conv2d_4_filter_read_block = 2;
  assign cparam_conv2d_4_filter_read_step = 16;
  assign cparam_conv2d_4_out_offset_values_0 = 0;
  assign cparam_conv2d_4_out_col_step = 64;
  assign cparam_conv2d_4_out_row_step = 1792;
  assign cparam_conv2d_4_out_bat_step = 50176;
  assign cparam_conv2d_4_out_och_step = 16;
  assign cparam_conv2d_4_out_write_size = 8;
  assign cparam_conv2d_4_out_write_size_res = 8;
  assign cparam_conv2d_4_out_write_block = 0;
  assign cparam_conv2d_4_keep_filter = 0;
  assign cparam_conv2d_4_keep_input = 1;
  assign cparam_conv2d_4_data_stationary = 0;
  assign cparam_conv2d_4_stream_num_ops = 8;
  assign cparam_conv2d_4_stream_num_ops_res = 8;
  assign cparam_conv2d_4_stream_num_ops_par = 8;
  assign cparam_conv2d_4_stream_num_ops_res_par = 8;
  assign cparam_conv2d_4_stream_reduce_size = 1;
  assign cparam_conv2d_4_stream_aligned_reduce_size = 2;
  assign cparam_conv2d_4_stream_omit_mask = 0;
  assign cparam_conv2d_4_col_select_initval = 2;
  assign cparam_conv2d_4_stride_col_par_col = 1;
  assign cparam_conv2d_4_stride_row_par_row = 1;
  assign cparam_conv2d_4_stride_col_mod_filter_num = 1;
  assign cparam_conv2d_4_filter_num_col_minus_stride_col_mod = 2;
  assign cparam_conv2d_4_inc_act_laddr_conds_0 = 1;
  assign cparam_conv2d_4_inc_act_laddr_conds_1 = 0;
  assign cparam_conv2d_4_inc_act_laddr_conds_2 = 0;
  assign cparam_conv2d_4_inc_act_laddr_conds_3 = 0;
  assign cparam_conv2d_4_inc_act_laddr_conds_4 = 1;
  assign cparam_conv2d_4_inc_act_laddr_conds_5 = 0;
  assign cparam_conv2d_4_inc_act_laddr_conds_6 = 0;
  assign cparam_conv2d_4_inc_act_laddr_conds_7 = 0;
  assign cparam_conv2d_4_inc_act_laddr_conds_8 = 1;
  assign cparam_conv2d_4_inc_act_laddr_conds_9 = 1;
  assign cparam_conv2d_4_inc_act_laddr_conds_10 = 0;
  assign cparam_conv2d_4_inc_act_laddr_conds_11 = 0;
  assign cparam_conv2d_4_inc_act_laddr_conds_12 = 0;
  assign cparam_conv2d_4_inc_act_laddr_conds_13 = 1;
  assign cparam_conv2d_4_inc_act_laddr_conds_14 = 0;
  assign cparam_conv2d_4_inc_act_laddr_conds_15 = 0;
  assign cparam_conv2d_4_inc_act_laddr_conds_16 = 0;
  assign cparam_conv2d_4_inc_act_laddr_conds_17 = 1;
  assign cparam_conv2d_4_inc_act_laddr_conds_18 = 1;
  assign cparam_conv2d_4_inc_act_laddr_conds_19 = 0;
  assign cparam_conv2d_4_inc_act_laddr_conds_20 = 0;
  assign cparam_conv2d_4_inc_act_laddr_conds_21 = 0;
  assign cparam_conv2d_4_inc_act_laddr_conds_22 = 1;
  assign cparam_conv2d_4_inc_act_laddr_conds_23 = 0;
  assign cparam_conv2d_4_inc_act_laddr_conds_24 = 0;
  assign cparam_conv2d_4_inc_act_laddr_conds_25 = 0;
  assign cparam_conv2d_4_inc_act_laddr_conds_26 = 1;
  assign cparam_conv2d_4_inc_act_laddr_small = 0;
  assign cparam_conv2d_4_inc_act_laddr_large = 2;
  assign cparam_conv2d_4_inc_out_laddr_col = 32;
  assign cparam_conv2d_4_stream_act_local_small_offset = 0;
  assign cparam_conv2d_4_stream_act_local_large_offset = -2;
  assign cparam_conv2d_4_stream_act_local_small_flags_0 = 0;
  assign cparam_conv2d_4_stream_act_local_small_flags_1 = 0;
  assign cparam_conv2d_4_stream_act_local_small_flags_2 = 1;
  assign cparam_conv2d_4_stream_act_local_large_flags_0 = 0;
  assign cparam_conv2d_4_stream_act_local_large_flags_1 = 0;
  assign cparam_conv2d_4_stream_act_local_large_flags_2 = 1;
  assign cparam_conv2d_4_inc_sync_out = 1;
  assign cparam_conv2d_4_inc_sync_out_res = 0;
  wire [5-1:0] cparam_max_pool_serial_6_act_num_col;
  wire [5-1:0] cparam_max_pool_serial_6_act_num_row;
  wire [2-1:0] cparam_max_pool_serial_6_stride_col;
  wire [2-1:0] cparam_max_pool_serial_6_stride_row;
  wire [4-1:0] cparam_max_pool_serial_6_out_num_col;
  wire [4-1:0] cparam_max_pool_serial_6_out_num_row;
  wire [1-1:0] cparam_max_pool_serial_6_pad_col_left;
  wire [1-1:0] cparam_max_pool_serial_6_pad_row_top;
  wire [5-1:0] cparam_max_pool_serial_6_max_col_count;
  wire [5-1:0] cparam_max_pool_serial_6_max_row_count;
  wire [1-1:0] cparam_max_pool_serial_6_max_bat_count;
  wire signed [32-1:0] cparam_max_pool_serial_6_act_offset_values_0;
  wire signed [32-1:0] cparam_max_pool_serial_6_act_offset_values_1;
  wire [12-1:0] cparam_max_pool_serial_6_act_row_step;
  wire [16-1:0] cparam_max_pool_serial_6_act_bat_step;
  wire [10-1:0] cparam_max_pool_serial_6_act_read_size;
  wire [6-1:0] cparam_max_pool_serial_6_act_read_block;
  wire [10-1:0] cparam_max_pool_serial_6_out_row_step;
  wire [14-1:0] cparam_max_pool_serial_6_out_bat_step;
  wire [9-1:0] cparam_max_pool_serial_6_out_write_size;
  wire [6-1:0] cparam_max_pool_serial_6_stream_size;
  wire [1-1:0] cparam_max_pool_serial_6_col_select_initval;
  wire [1-1:0] cparam_max_pool_serial_6_stride_col_mod_ksize;
  wire [2-1:0] cparam_max_pool_serial_6_ksize_col_minus_stride_col_mod;
  wire [1-1:0] cparam_max_pool_serial_6_local_pad_offset;
  wire [7-1:0] cparam_max_pool_serial_6_inc_act_laddr;
  wire [6-1:0] cparam_max_pool_serial_6_inc_out_laddr;
  assign cparam_max_pool_serial_6_act_num_col = 28;
  assign cparam_max_pool_serial_6_act_num_row = 28;
  assign cparam_max_pool_serial_6_stride_col = 2;
  assign cparam_max_pool_serial_6_stride_row = 2;
  assign cparam_max_pool_serial_6_out_num_col = 14;
  assign cparam_max_pool_serial_6_out_num_row = 14;
  assign cparam_max_pool_serial_6_pad_col_left = 0;
  assign cparam_max_pool_serial_6_pad_row_top = 0;
  assign cparam_max_pool_serial_6_max_col_count = 25;
  assign cparam_max_pool_serial_6_max_row_count = 25;
  assign cparam_max_pool_serial_6_max_bat_count = 0;
  assign cparam_max_pool_serial_6_act_offset_values_0 = 0;
  assign cparam_max_pool_serial_6_act_offset_values_1 = 1792;
  assign cparam_max_pool_serial_6_act_row_step = 3584;
  assign cparam_max_pool_serial_6_act_bat_step = 50176;
  assign cparam_max_pool_serial_6_act_read_size = 896;
  assign cparam_max_pool_serial_6_act_read_block = 32;
  assign cparam_max_pool_serial_6_out_row_step = 896;
  assign cparam_max_pool_serial_6_out_bat_step = 12544;
  assign cparam_max_pool_serial_6_out_write_size = 448;
  assign cparam_max_pool_serial_6_stream_size = 32;
  assign cparam_max_pool_serial_6_col_select_initval = 0;
  assign cparam_max_pool_serial_6_stride_col_mod_ksize = 0;
  assign cparam_max_pool_serial_6_ksize_col_minus_stride_col_mod = 2;
  assign cparam_max_pool_serial_6_local_pad_offset = 0;
  assign cparam_max_pool_serial_6_inc_act_laddr = 64;
  assign cparam_max_pool_serial_6_inc_out_laddr = 32;
  wire [1-1:0] cparam_matmul_11_act_num_col;
  wire [1-1:0] cparam_matmul_11_act_num_row;
  wire [8-1:0] cparam_matmul_11_filter_num_och;
  wire [1-1:0] cparam_matmul_11_bias_scala;
  wire [8-1:0] cparam_matmul_11_bias_num;
  wire [1-1:0] cparam_matmul_11_scale_scala;
  wire [8-1:0] cparam_matmul_11_scale_num;
  wire [1-1:0] cparam_matmul_11_vshamt_mul_scala;
  wire [1-1:0] cparam_matmul_11_vshamt_mul_num;
  wire [1-1:0] cparam_matmul_11_vshamt_sum_scala;
  wire [1-1:0] cparam_matmul_11_vshamt_sum_num;
  wire [1-1:0] cparam_matmul_11_vshamt_out_scala;
  wire [1-1:0] cparam_matmul_11_vshamt_out_num;
  wire [1-1:0] cparam_matmul_11_cshamt_mul_value;
  wire [1-1:0] cparam_matmul_11_cshamt_sum_value;
  wire [5-1:0] cparam_matmul_11_cshamt_out_value;
  wire [1-1:0] cparam_matmul_11_act_func_index;
  wire [1-1:0] cparam_matmul_11_out_num_col;
  wire [1-1:0] cparam_matmul_11_out_num_row;
  wire [1-1:0] cparam_matmul_11_pad_col_left;
  wire [1-1:0] cparam_matmul_11_pad_row_top;
  wire [1-1:0] cparam_matmul_11_max_col_count;
  wire [1-1:0] cparam_matmul_11_max_row_count;
  wire [1-1:0] cparam_matmul_11_max_bat_count;
  wire [7-1:0] cparam_matmul_11_max_och_count;
  wire [8-1:0] cparam_matmul_11_och_count_step;
  wire [1-1:0] cparam_matmul_11_dma_flag_conds_0;
  wire signed [32-1:0] cparam_matmul_11_act_offset_values_0;
  wire [14-1:0] cparam_matmul_11_act_row_step;
  wire [14-1:0] cparam_matmul_11_act_bat_step;
  wire [13-1:0] cparam_matmul_11_act_read_size;
  wire [13-1:0] cparam_matmul_11_act_read_block;
  wire [13-1:0] cparam_matmul_11_act_read_step;
  wire [15-1:0] cparam_matmul_11_filter_base_step;
  wire [14-1:0] cparam_matmul_11_filter_read_size;
  wire [13-1:0] cparam_matmul_11_filter_read_block;
  wire [14-1:0] cparam_matmul_11_filter_read_step;
  wire [1-1:0] cparam_matmul_11_out_offset_values_0;
  wire [9-1:0] cparam_matmul_11_out_col_step;
  wire [9-1:0] cparam_matmul_11_out_row_step;
  wire [9-1:0] cparam_matmul_11_out_bat_step;
  wire [5-1:0] cparam_matmul_11_out_och_step;
  wire [4-1:0] cparam_matmul_11_out_write_size;
  wire [4-1:0] cparam_matmul_11_out_write_size_res;
  wire [4-1:0] cparam_matmul_11_out_write_block;
  wire [1-1:0] cparam_matmul_11_keep_filter;
  wire [1-1:0] cparam_matmul_11_keep_input;
  wire [1-1:0] cparam_matmul_11_data_stationary;
  wire [4-1:0] cparam_matmul_11_stream_num_ops;
  wire [4-1:0] cparam_matmul_11_stream_num_ops_res;
  wire [4-1:0] cparam_matmul_11_stream_num_ops_par;
  wire [4-1:0] cparam_matmul_11_stream_num_ops_res_par;
  wire [13-1:0] cparam_matmul_11_stream_reduce_size;
  wire [13-1:0] cparam_matmul_11_stream_aligned_reduce_size;
  wire [1-1:0] cparam_matmul_11_stream_omit_mask;
  wire [1-1:0] cparam_matmul_11_col_select_initval;
  wire [1-1:0] cparam_matmul_11_stride_col_par_col;
  wire [1-1:0] cparam_matmul_11_stride_row_par_row;
  wire [1-1:0] cparam_matmul_11_stride_col_mod_filter_num;
  wire [1-1:0] cparam_matmul_11_filter_num_col_minus_stride_col_mod;
  wire [1-1:0] cparam_matmul_11_inc_act_laddr_conds_0;
  wire [13-1:0] cparam_matmul_11_inc_act_laddr_small;
  wire [13-1:0] cparam_matmul_11_inc_act_laddr_large;
  wire [8-1:0] cparam_matmul_11_inc_out_laddr_col;
  wire [1-1:0] cparam_matmul_11_stream_act_local_small_offset;
  wire [1-1:0] cparam_matmul_11_stream_act_local_large_offset;
  wire [1-1:0] cparam_matmul_11_stream_act_local_small_flags_0;
  wire [1-1:0] cparam_matmul_11_stream_act_local_large_flags_0;
  wire [1-1:0] cparam_matmul_11_inc_sync_out;
  wire [1-1:0] cparam_matmul_11_inc_sync_out_res;
  reg [1-1:0] matmul_11_control_param_index;
  assign cparam_matmul_11_act_num_col = (matmul_11_control_param_index == 0)? 32'h1 : 32'h1;
  assign cparam_matmul_11_act_num_row = (matmul_11_control_param_index == 0)? 32'h1 : 32'h1;
  assign cparam_matmul_11_filter_num_och = (matmul_11_control_param_index == 0)? 32'h80 : 32'ha;
  assign cparam_matmul_11_bias_scala = (matmul_11_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_11_bias_num = (matmul_11_control_param_index == 0)? 32'h80 : 32'ha;
  assign cparam_matmul_11_scale_scala = (matmul_11_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_11_scale_num = (matmul_11_control_param_index == 0)? 32'h80 : 32'ha;
  assign cparam_matmul_11_vshamt_mul_scala = (matmul_11_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_11_vshamt_mul_num = (matmul_11_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_11_vshamt_sum_scala = (matmul_11_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_11_vshamt_sum_num = (matmul_11_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_11_vshamt_out_scala = (matmul_11_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_11_vshamt_out_num = (matmul_11_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_11_cshamt_mul_value = (matmul_11_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_11_cshamt_sum_value = (matmul_11_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_11_cshamt_out_value = (matmul_11_control_param_index == 0)? 32'h1d : 32'h1d;
  assign cparam_matmul_11_act_func_index = (matmul_11_control_param_index == 0)? 32'h0 : 32'h1;
  assign cparam_matmul_11_out_num_col = (matmul_11_control_param_index == 0)? 32'h1 : 32'h1;
  assign cparam_matmul_11_out_num_row = (matmul_11_control_param_index == 0)? 32'h1 : 32'h1;
  assign cparam_matmul_11_pad_col_left = (matmul_11_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_11_pad_row_top = (matmul_11_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_11_max_col_count = (matmul_11_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_11_max_row_count = (matmul_11_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_11_max_bat_count = (matmul_11_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_11_max_och_count = (matmul_11_control_param_index == 0)? 32'h7e : 32'h0;
  assign cparam_matmul_11_och_count_step = (matmul_11_control_param_index == 0)? 32'h2 : 32'h80;
  assign cparam_matmul_11_dma_flag_conds_0 = (matmul_11_control_param_index == 0)? 32'h1 : 32'h1;
  assign cparam_matmul_11_act_offset_values_0 = (matmul_11_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_11_act_row_step = (matmul_11_control_param_index == 0)? 32'h3100 : 32'h100;
  assign cparam_matmul_11_act_bat_step = (matmul_11_control_param_index == 0)? 32'h3100 : 32'h100;
  assign cparam_matmul_11_act_read_size = (matmul_11_control_param_index == 0)? 32'h1880 : 32'h80;
  assign cparam_matmul_11_act_read_block = (matmul_11_control_param_index == 0)? 32'h1880 : 32'h80;
  assign cparam_matmul_11_act_read_step = (matmul_11_control_param_index == 0)? 32'h1880 : 32'h80;
  assign cparam_matmul_11_filter_base_step = (matmul_11_control_param_index == 0)? 32'h6200 : 32'ha00;
  assign cparam_matmul_11_filter_read_size = (matmul_11_control_param_index == 0)? 32'h3100 : 32'h500;
  assign cparam_matmul_11_filter_read_block = (matmul_11_control_param_index == 0)? 32'h1880 : 32'h80;
  assign cparam_matmul_11_filter_read_step = (matmul_11_control_param_index == 0)? 32'h3100 : 32'h500;
  assign cparam_matmul_11_out_offset_values_0 = (matmul_11_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_11_out_col_step = (matmul_11_control_param_index == 0)? 32'h100 : 32'h14;
  assign cparam_matmul_11_out_row_step = (matmul_11_control_param_index == 0)? 32'h100 : 32'h14;
  assign cparam_matmul_11_out_bat_step = (matmul_11_control_param_index == 0)? 32'h100 : 32'h14;
  assign cparam_matmul_11_out_och_step = (matmul_11_control_param_index == 0)? 32'h4 : 32'h14;
  assign cparam_matmul_11_out_write_size = (matmul_11_control_param_index == 0)? 32'h2 : 32'ha;
  assign cparam_matmul_11_out_write_size_res = (matmul_11_control_param_index == 0)? 32'h2 : 32'ha;
  assign cparam_matmul_11_out_write_block = (matmul_11_control_param_index == 0)? 32'h0 : 32'ha;
  assign cparam_matmul_11_keep_filter = (matmul_11_control_param_index == 0)? 32'h0 : 32'h1;
  assign cparam_matmul_11_keep_input = (matmul_11_control_param_index == 0)? 32'h1 : 32'h1;
  assign cparam_matmul_11_data_stationary = (matmul_11_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_11_stream_num_ops = (matmul_11_control_param_index == 0)? 32'h2 : 32'ha;
  assign cparam_matmul_11_stream_num_ops_res = (matmul_11_control_param_index == 0)? 32'h2 : 32'ha;
  assign cparam_matmul_11_stream_num_ops_par = (matmul_11_control_param_index == 0)? 32'h2 : 32'ha;
  assign cparam_matmul_11_stream_num_ops_res_par = (matmul_11_control_param_index == 0)? 32'h2 : 32'ha;
  assign cparam_matmul_11_stream_reduce_size = (matmul_11_control_param_index == 0)? 32'h1880 : 32'h80;
  assign cparam_matmul_11_stream_aligned_reduce_size = (matmul_11_control_param_index == 0)? 32'h1880 : 32'h80;
  assign cparam_matmul_11_stream_omit_mask = (matmul_11_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_11_col_select_initval = (matmul_11_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_11_stride_col_par_col = (matmul_11_control_param_index == 0)? 32'h1 : 32'h1;
  assign cparam_matmul_11_stride_row_par_row = (matmul_11_control_param_index == 0)? 32'h1 : 32'h1;
  assign cparam_matmul_11_stride_col_mod_filter_num = (matmul_11_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_11_filter_num_col_minus_stride_col_mod = (matmul_11_control_param_index == 0)? 32'h1 : 32'h1;
  assign cparam_matmul_11_inc_act_laddr_conds_0 = (matmul_11_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_11_inc_act_laddr_small = (matmul_11_control_param_index == 0)? 32'h1880 : 32'h80;
  assign cparam_matmul_11_inc_act_laddr_large = (matmul_11_control_param_index == 0)? 32'h1880 : 32'h80;
  assign cparam_matmul_11_inc_out_laddr_col = (matmul_11_control_param_index == 0)? 32'h80 : 32'ha;
  assign cparam_matmul_11_stream_act_local_small_offset = (matmul_11_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_11_stream_act_local_large_offset = (matmul_11_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_11_stream_act_local_small_flags_0 = (matmul_11_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_11_stream_act_local_large_flags_0 = (matmul_11_control_param_index == 0)? 32'h0 : 32'h0;
  assign cparam_matmul_11_inc_sync_out = (matmul_11_control_param_index == 0)? 32'h1 : 32'h1;
  assign cparam_matmul_11_inc_sync_out_res = (matmul_11_control_param_index == 0)? 32'h0 : 32'h0;
  reg _acc_14_stream_ivalid;
  wire _acc_14_stream_oready;
  wire _acc_14_stream_internal_oready;
  assign _acc_14_stream_internal_oready = 1;
  reg [32-1:0] _acc_14_fsm;
  localparam _acc_14_fsm_init = 0;
  wire _acc_14_run_flag;
  assign _acc_14_run_flag = 0;
  reg _acc_14_source_start;
  wire _acc_14_source_stop;
  reg _acc_14_source_busy;
  wire _acc_14_sink_start;
  wire _acc_14_sink_stop;
  wire _acc_14_sink_busy;
  wire _acc_14_busy;
  reg _acc_14_busy_reg;
  wire _acc_14_is_root;
  reg _acc_14_x_idle;
  reg [33-1:0] _acc_14_x_source_count;
  reg [5-1:0] _acc_14_x_source_mode;
  reg [16-1:0] _acc_14_x_source_generator_id;
  reg [32-1:0] _acc_14_x_source_offset;
  reg [33-1:0] _acc_14_x_source_size;
  reg [32-1:0] _acc_14_x_source_stride;
  reg [32-1:0] _acc_14_x_source_offset_buf;
  reg [33-1:0] _acc_14_x_source_size_buf;
  reg [32-1:0] _acc_14_x_source_stride_buf;
  reg [8-1:0] _acc_14_x_source_sel;
  reg [32-1:0] _acc_14_x_source_ram_raddr;
  reg _acc_14_x_source_ram_renable;
  wire [64-1:0] _acc_14_x_source_ram_rdata;
  reg _acc_14_x_source_fifo_deq;
  wire [64-1:0] _acc_14_x_source_fifo_rdata;
  reg [64-1:0] _acc_14_x_source_empty_data;
  reg _acc_14_rshift_idle;
  reg [33-1:0] _acc_14_rshift_source_count;
  reg [5-1:0] _acc_14_rshift_source_mode;
  reg [16-1:0] _acc_14_rshift_source_generator_id;
  reg [32-1:0] _acc_14_rshift_source_offset;
  reg [33-1:0] _acc_14_rshift_source_size;
  reg [32-1:0] _acc_14_rshift_source_stride;
  reg [32-1:0] _acc_14_rshift_source_offset_buf;
  reg [33-1:0] _acc_14_rshift_source_size_buf;
  reg [32-1:0] _acc_14_rshift_source_stride_buf;
  reg [8-1:0] _acc_14_rshift_source_sel;
  reg [32-1:0] _acc_14_rshift_source_ram_raddr;
  reg _acc_14_rshift_source_ram_renable;
  wire [32-1:0] _acc_14_rshift_source_ram_rdata;
  reg _acc_14_rshift_source_fifo_deq;
  wire [32-1:0] _acc_14_rshift_source_fifo_rdata;
  reg [32-1:0] _acc_14_rshift_source_empty_data;
  reg [32-1:0] _acc_14_size_next_parameter_data;
  reg [33-1:0] _acc_14_sum_sink_count;
  reg [5-1:0] _acc_14_sum_sink_mode;
  reg [16-1:0] _acc_14_sum_sink_generator_id;
  reg [32-1:0] _acc_14_sum_sink_offset;
  reg [33-1:0] _acc_14_sum_sink_size;
  reg [32-1:0] _acc_14_sum_sink_stride;
  reg [32-1:0] _acc_14_sum_sink_offset_buf;
  reg [33-1:0] _acc_14_sum_sink_size_buf;
  reg [32-1:0] _acc_14_sum_sink_stride_buf;
  reg [8-1:0] _acc_14_sum_sink_sel;
  reg [32-1:0] _acc_14_sum_sink_waddr;
  reg _acc_14_sum_sink_wenable;
  reg [64-1:0] _acc_14_sum_sink_wdata;
  reg _acc_14_sum_sink_fifo_enq;
  reg [64-1:0] _acc_14_sum_sink_fifo_wdata;
  reg [64-1:0] _acc_14_sum_sink_immediate;
  reg [33-1:0] _acc_14_valid_sink_count;
  reg [5-1:0] _acc_14_valid_sink_mode;
  reg [16-1:0] _acc_14_valid_sink_generator_id;
  reg [32-1:0] _acc_14_valid_sink_offset;
  reg [33-1:0] _acc_14_valid_sink_size;
  reg [32-1:0] _acc_14_valid_sink_stride;
  reg [32-1:0] _acc_14_valid_sink_offset_buf;
  reg [33-1:0] _acc_14_valid_sink_size_buf;
  reg [32-1:0] _acc_14_valid_sink_stride_buf;
  reg [8-1:0] _acc_14_valid_sink_sel;
  reg [32-1:0] _acc_14_valid_sink_waddr;
  reg _acc_14_valid_sink_wenable;
  reg [1-1:0] _acc_14_valid_sink_wdata;
  reg _acc_14_valid_sink_fifo_enq;
  reg [1-1:0] _acc_14_valid_sink_fifo_wdata;
  reg [1-1:0] _acc_14_valid_sink_immediate;
  reg _add_tree_15_stream_ivalid;
  wire _add_tree_15_stream_oready;
  wire _add_tree_15_stream_internal_oready;
  assign _add_tree_15_stream_internal_oready = 1;
  reg [32-1:0] _add_tree_15_fsm;
  localparam _add_tree_15_fsm_init = 0;
  wire _add_tree_15_run_flag;
  assign _add_tree_15_run_flag = 0;
  reg _add_tree_15_source_start;
  wire _add_tree_15_source_stop;
  reg _add_tree_15_source_busy;
  wire _add_tree_15_sink_start;
  wire _add_tree_15_sink_stop;
  wire _add_tree_15_sink_busy;
  wire _add_tree_15_busy;
  reg _add_tree_15_busy_reg;
  wire _add_tree_15_is_root;
  reg _add_tree_15_var0_idle;
  reg [33-1:0] _add_tree_15_var0_source_count;
  reg [5-1:0] _add_tree_15_var0_source_mode;
  reg [16-1:0] _add_tree_15_var0_source_generator_id;
  reg [32-1:0] _add_tree_15_var0_source_offset;
  reg [33-1:0] _add_tree_15_var0_source_size;
  reg [32-1:0] _add_tree_15_var0_source_stride;
  reg [32-1:0] _add_tree_15_var0_source_offset_buf;
  reg [33-1:0] _add_tree_15_var0_source_size_buf;
  reg [32-1:0] _add_tree_15_var0_source_stride_buf;
  reg [8-1:0] _add_tree_15_var0_source_sel;
  reg [32-1:0] _add_tree_15_var0_source_ram_raddr;
  reg _add_tree_15_var0_source_ram_renable;
  wire [64-1:0] _add_tree_15_var0_source_ram_rdata;
  reg _add_tree_15_var0_source_fifo_deq;
  wire [64-1:0] _add_tree_15_var0_source_fifo_rdata;
  reg [64-1:0] _add_tree_15_var0_source_empty_data;
  reg [33-1:0] _add_tree_15_sum_sink_count;
  reg [5-1:0] _add_tree_15_sum_sink_mode;
  reg [16-1:0] _add_tree_15_sum_sink_generator_id;
  reg [32-1:0] _add_tree_15_sum_sink_offset;
  reg [33-1:0] _add_tree_15_sum_sink_size;
  reg [32-1:0] _add_tree_15_sum_sink_stride;
  reg [32-1:0] _add_tree_15_sum_sink_offset_buf;
  reg [33-1:0] _add_tree_15_sum_sink_size_buf;
  reg [32-1:0] _add_tree_15_sum_sink_stride_buf;
  reg [8-1:0] _add_tree_15_sum_sink_sel;
  reg [32-1:0] _add_tree_15_sum_sink_waddr;
  reg _add_tree_15_sum_sink_wenable;
  reg [64-1:0] _add_tree_15_sum_sink_wdata;
  reg _add_tree_15_sum_sink_fifo_enq;
  reg [64-1:0] _add_tree_15_sum_sink_fifo_wdata;
  reg [64-1:0] _add_tree_15_sum_sink_immediate;
  reg _add_tree_16_stream_ivalid;
  wire _add_tree_16_stream_oready;
  wire _add_tree_16_stream_internal_oready;
  assign _add_tree_16_stream_internal_oready = 1;
  reg [32-1:0] _add_tree_16_fsm;
  localparam _add_tree_16_fsm_init = 0;
  wire _add_tree_16_run_flag;
  assign _add_tree_16_run_flag = 0;
  reg _add_tree_16_source_start;
  wire _add_tree_16_source_stop;
  reg _add_tree_16_source_busy;
  wire _add_tree_16_sink_start;
  wire _add_tree_16_sink_stop;
  wire _add_tree_16_sink_busy;
  wire _add_tree_16_busy;
  reg _add_tree_16_busy_reg;
  wire _add_tree_16_is_root;
  reg _add_tree_16_var0_idle;
  reg [33-1:0] _add_tree_16_var0_source_count;
  reg [5-1:0] _add_tree_16_var0_source_mode;
  reg [16-1:0] _add_tree_16_var0_source_generator_id;
  reg [32-1:0] _add_tree_16_var0_source_offset;
  reg [33-1:0] _add_tree_16_var0_source_size;
  reg [32-1:0] _add_tree_16_var0_source_stride;
  reg [32-1:0] _add_tree_16_var0_source_offset_buf;
  reg [33-1:0] _add_tree_16_var0_source_size_buf;
  reg [32-1:0] _add_tree_16_var0_source_stride_buf;
  reg [8-1:0] _add_tree_16_var0_source_sel;
  reg [32-1:0] _add_tree_16_var0_source_ram_raddr;
  reg _add_tree_16_var0_source_ram_renable;
  wire [64-1:0] _add_tree_16_var0_source_ram_rdata;
  reg _add_tree_16_var0_source_fifo_deq;
  wire [64-1:0] _add_tree_16_var0_source_fifo_rdata;
  reg [64-1:0] _add_tree_16_var0_source_empty_data;
  reg _add_tree_16_var1_idle;
  reg [33-1:0] _add_tree_16_var1_source_count;
  reg [5-1:0] _add_tree_16_var1_source_mode;
  reg [16-1:0] _add_tree_16_var1_source_generator_id;
  reg [32-1:0] _add_tree_16_var1_source_offset;
  reg [33-1:0] _add_tree_16_var1_source_size;
  reg [32-1:0] _add_tree_16_var1_source_stride;
  reg [32-1:0] _add_tree_16_var1_source_offset_buf;
  reg [33-1:0] _add_tree_16_var1_source_size_buf;
  reg [32-1:0] _add_tree_16_var1_source_stride_buf;
  reg [8-1:0] _add_tree_16_var1_source_sel;
  reg [32-1:0] _add_tree_16_var1_source_ram_raddr;
  reg _add_tree_16_var1_source_ram_renable;
  wire [64-1:0] _add_tree_16_var1_source_ram_rdata;
  reg _add_tree_16_var1_source_fifo_deq;
  wire [64-1:0] _add_tree_16_var1_source_fifo_rdata;
  reg [64-1:0] _add_tree_16_var1_source_empty_data;
  reg _add_tree_16_var2_idle;
  reg [33-1:0] _add_tree_16_var2_source_count;
  reg [5-1:0] _add_tree_16_var2_source_mode;
  reg [16-1:0] _add_tree_16_var2_source_generator_id;
  reg [32-1:0] _add_tree_16_var2_source_offset;
  reg [33-1:0] _add_tree_16_var2_source_size;
  reg [32-1:0] _add_tree_16_var2_source_stride;
  reg [32-1:0] _add_tree_16_var2_source_offset_buf;
  reg [33-1:0] _add_tree_16_var2_source_size_buf;
  reg [32-1:0] _add_tree_16_var2_source_stride_buf;
  reg [8-1:0] _add_tree_16_var2_source_sel;
  reg [32-1:0] _add_tree_16_var2_source_ram_raddr;
  reg _add_tree_16_var2_source_ram_renable;
  wire [64-1:0] _add_tree_16_var2_source_ram_rdata;
  reg _add_tree_16_var2_source_fifo_deq;
  wire [64-1:0] _add_tree_16_var2_source_fifo_rdata;
  reg [64-1:0] _add_tree_16_var2_source_empty_data;
  reg _add_tree_16_var3_idle;
  reg [33-1:0] _add_tree_16_var3_source_count;
  reg [5-1:0] _add_tree_16_var3_source_mode;
  reg [16-1:0] _add_tree_16_var3_source_generator_id;
  reg [32-1:0] _add_tree_16_var3_source_offset;
  reg [33-1:0] _add_tree_16_var3_source_size;
  reg [32-1:0] _add_tree_16_var3_source_stride;
  reg [32-1:0] _add_tree_16_var3_source_offset_buf;
  reg [33-1:0] _add_tree_16_var3_source_size_buf;
  reg [32-1:0] _add_tree_16_var3_source_stride_buf;
  reg [8-1:0] _add_tree_16_var3_source_sel;
  reg [32-1:0] _add_tree_16_var3_source_ram_raddr;
  reg _add_tree_16_var3_source_ram_renable;
  wire [64-1:0] _add_tree_16_var3_source_ram_rdata;
  reg _add_tree_16_var3_source_fifo_deq;
  wire [64-1:0] _add_tree_16_var3_source_fifo_rdata;
  reg [64-1:0] _add_tree_16_var3_source_empty_data;
  reg _add_tree_16_var4_idle;
  reg [33-1:0] _add_tree_16_var4_source_count;
  reg [5-1:0] _add_tree_16_var4_source_mode;
  reg [16-1:0] _add_tree_16_var4_source_generator_id;
  reg [32-1:0] _add_tree_16_var4_source_offset;
  reg [33-1:0] _add_tree_16_var4_source_size;
  reg [32-1:0] _add_tree_16_var4_source_stride;
  reg [32-1:0] _add_tree_16_var4_source_offset_buf;
  reg [33-1:0] _add_tree_16_var4_source_size_buf;
  reg [32-1:0] _add_tree_16_var4_source_stride_buf;
  reg [8-1:0] _add_tree_16_var4_source_sel;
  reg [32-1:0] _add_tree_16_var4_source_ram_raddr;
  reg _add_tree_16_var4_source_ram_renable;
  wire [64-1:0] _add_tree_16_var4_source_ram_rdata;
  reg _add_tree_16_var4_source_fifo_deq;
  wire [64-1:0] _add_tree_16_var4_source_fifo_rdata;
  reg [64-1:0] _add_tree_16_var4_source_empty_data;
  reg _add_tree_16_var5_idle;
  reg [33-1:0] _add_tree_16_var5_source_count;
  reg [5-1:0] _add_tree_16_var5_source_mode;
  reg [16-1:0] _add_tree_16_var5_source_generator_id;
  reg [32-1:0] _add_tree_16_var5_source_offset;
  reg [33-1:0] _add_tree_16_var5_source_size;
  reg [32-1:0] _add_tree_16_var5_source_stride;
  reg [32-1:0] _add_tree_16_var5_source_offset_buf;
  reg [33-1:0] _add_tree_16_var5_source_size_buf;
  reg [32-1:0] _add_tree_16_var5_source_stride_buf;
  reg [8-1:0] _add_tree_16_var5_source_sel;
  reg [32-1:0] _add_tree_16_var5_source_ram_raddr;
  reg _add_tree_16_var5_source_ram_renable;
  wire [64-1:0] _add_tree_16_var5_source_ram_rdata;
  reg _add_tree_16_var5_source_fifo_deq;
  wire [64-1:0] _add_tree_16_var5_source_fifo_rdata;
  reg [64-1:0] _add_tree_16_var5_source_empty_data;
  reg _add_tree_16_var6_idle;
  reg [33-1:0] _add_tree_16_var6_source_count;
  reg [5-1:0] _add_tree_16_var6_source_mode;
  reg [16-1:0] _add_tree_16_var6_source_generator_id;
  reg [32-1:0] _add_tree_16_var6_source_offset;
  reg [33-1:0] _add_tree_16_var6_source_size;
  reg [32-1:0] _add_tree_16_var6_source_stride;
  reg [32-1:0] _add_tree_16_var6_source_offset_buf;
  reg [33-1:0] _add_tree_16_var6_source_size_buf;
  reg [32-1:0] _add_tree_16_var6_source_stride_buf;
  reg [8-1:0] _add_tree_16_var6_source_sel;
  reg [32-1:0] _add_tree_16_var6_source_ram_raddr;
  reg _add_tree_16_var6_source_ram_renable;
  wire [64-1:0] _add_tree_16_var6_source_ram_rdata;
  reg _add_tree_16_var6_source_fifo_deq;
  wire [64-1:0] _add_tree_16_var6_source_fifo_rdata;
  reg [64-1:0] _add_tree_16_var6_source_empty_data;
  reg _add_tree_16_var7_idle;
  reg [33-1:0] _add_tree_16_var7_source_count;
  reg [5-1:0] _add_tree_16_var7_source_mode;
  reg [16-1:0] _add_tree_16_var7_source_generator_id;
  reg [32-1:0] _add_tree_16_var7_source_offset;
  reg [33-1:0] _add_tree_16_var7_source_size;
  reg [32-1:0] _add_tree_16_var7_source_stride;
  reg [32-1:0] _add_tree_16_var7_source_offset_buf;
  reg [33-1:0] _add_tree_16_var7_source_size_buf;
  reg [32-1:0] _add_tree_16_var7_source_stride_buf;
  reg [8-1:0] _add_tree_16_var7_source_sel;
  reg [32-1:0] _add_tree_16_var7_source_ram_raddr;
  reg _add_tree_16_var7_source_ram_renable;
  wire [64-1:0] _add_tree_16_var7_source_ram_rdata;
  reg _add_tree_16_var7_source_fifo_deq;
  wire [64-1:0] _add_tree_16_var7_source_fifo_rdata;
  reg [64-1:0] _add_tree_16_var7_source_empty_data;
  reg _add_tree_16_var8_idle;
  reg [33-1:0] _add_tree_16_var8_source_count;
  reg [5-1:0] _add_tree_16_var8_source_mode;
  reg [16-1:0] _add_tree_16_var8_source_generator_id;
  reg [32-1:0] _add_tree_16_var8_source_offset;
  reg [33-1:0] _add_tree_16_var8_source_size;
  reg [32-1:0] _add_tree_16_var8_source_stride;
  reg [32-1:0] _add_tree_16_var8_source_offset_buf;
  reg [33-1:0] _add_tree_16_var8_source_size_buf;
  reg [32-1:0] _add_tree_16_var8_source_stride_buf;
  reg [8-1:0] _add_tree_16_var8_source_sel;
  reg [32-1:0] _add_tree_16_var8_source_ram_raddr;
  reg _add_tree_16_var8_source_ram_renable;
  wire [64-1:0] _add_tree_16_var8_source_ram_rdata;
  reg _add_tree_16_var8_source_fifo_deq;
  wire [64-1:0] _add_tree_16_var8_source_fifo_rdata;
  reg [64-1:0] _add_tree_16_var8_source_empty_data;
  reg [33-1:0] _add_tree_16_sum_sink_count;
  reg [5-1:0] _add_tree_16_sum_sink_mode;
  reg [16-1:0] _add_tree_16_sum_sink_generator_id;
  reg [32-1:0] _add_tree_16_sum_sink_offset;
  reg [33-1:0] _add_tree_16_sum_sink_size;
  reg [32-1:0] _add_tree_16_sum_sink_stride;
  reg [32-1:0] _add_tree_16_sum_sink_offset_buf;
  reg [33-1:0] _add_tree_16_sum_sink_size_buf;
  reg [32-1:0] _add_tree_16_sum_sink_stride_buf;
  reg [8-1:0] _add_tree_16_sum_sink_sel;
  reg [32-1:0] _add_tree_16_sum_sink_waddr;
  reg _add_tree_16_sum_sink_wenable;
  reg [64-1:0] _add_tree_16_sum_sink_wdata;
  reg _add_tree_16_sum_sink_fifo_enq;
  reg [64-1:0] _add_tree_16_sum_sink_fifo_wdata;
  reg [64-1:0] _add_tree_16_sum_sink_immediate;
  reg _mul_rshift_round_clip_17_stream_ivalid;
  wire _mul_rshift_round_clip_17_stream_oready;
  wire _mul_rshift_round_clip_17_stream_internal_oready;
  assign _mul_rshift_round_clip_17_stream_internal_oready = 1;
  reg [32-1:0] _mul_rshift_round_clip_17_fsm;
  localparam _mul_rshift_round_clip_17_fsm_init = 0;
  wire _mul_rshift_round_clip_17_run_flag;
  assign _mul_rshift_round_clip_17_run_flag = 0;
  reg _mul_rshift_round_clip_17_source_start;
  wire _mul_rshift_round_clip_17_source_stop;
  reg _mul_rshift_round_clip_17_source_busy;
  wire _mul_rshift_round_clip_17_sink_start;
  wire _mul_rshift_round_clip_17_sink_stop;
  wire _mul_rshift_round_clip_17_sink_busy;
  wire _mul_rshift_round_clip_17_busy;
  reg _mul_rshift_round_clip_17_busy_reg;
  wire _mul_rshift_round_clip_17_is_root;
  reg _mul_rshift_round_clip_17_x_idle;
  reg [33-1:0] _mul_rshift_round_clip_17_x_source_count;
  reg [5-1:0] _mul_rshift_round_clip_17_x_source_mode;
  reg [16-1:0] _mul_rshift_round_clip_17_x_source_generator_id;
  reg [32-1:0] _mul_rshift_round_clip_17_x_source_offset;
  reg [33-1:0] _mul_rshift_round_clip_17_x_source_size;
  reg [32-1:0] _mul_rshift_round_clip_17_x_source_stride;
  reg [32-1:0] _mul_rshift_round_clip_17_x_source_offset_buf;
  reg [33-1:0] _mul_rshift_round_clip_17_x_source_size_buf;
  reg [32-1:0] _mul_rshift_round_clip_17_x_source_stride_buf;
  reg [8-1:0] _mul_rshift_round_clip_17_x_source_sel;
  reg [32-1:0] _mul_rshift_round_clip_17_x_source_ram_raddr;
  reg _mul_rshift_round_clip_17_x_source_ram_renable;
  wire [64-1:0] _mul_rshift_round_clip_17_x_source_ram_rdata;
  reg _mul_rshift_round_clip_17_x_source_fifo_deq;
  wire [64-1:0] _mul_rshift_round_clip_17_x_source_fifo_rdata;
  reg [64-1:0] _mul_rshift_round_clip_17_x_source_empty_data;
  reg _mul_rshift_round_clip_17_y_idle;
  reg [33-1:0] _mul_rshift_round_clip_17_y_source_count;
  reg [5-1:0] _mul_rshift_round_clip_17_y_source_mode;
  reg [16-1:0] _mul_rshift_round_clip_17_y_source_generator_id;
  reg [32-1:0] _mul_rshift_round_clip_17_y_source_offset;
  reg [33-1:0] _mul_rshift_round_clip_17_y_source_size;
  reg [32-1:0] _mul_rshift_round_clip_17_y_source_stride;
  reg [32-1:0] _mul_rshift_round_clip_17_y_source_offset_buf;
  reg [33-1:0] _mul_rshift_round_clip_17_y_source_size_buf;
  reg [32-1:0] _mul_rshift_round_clip_17_y_source_stride_buf;
  reg [8-1:0] _mul_rshift_round_clip_17_y_source_sel;
  reg [32-1:0] _mul_rshift_round_clip_17_y_source_ram_raddr;
  reg _mul_rshift_round_clip_17_y_source_ram_renable;
  wire [16-1:0] _mul_rshift_round_clip_17_y_source_ram_rdata;
  reg _mul_rshift_round_clip_17_y_source_fifo_deq;
  wire [16-1:0] _mul_rshift_round_clip_17_y_source_fifo_rdata;
  reg [16-1:0] _mul_rshift_round_clip_17_y_source_empty_data;
  reg _mul_rshift_round_clip_17_rshift_idle;
  reg [33-1:0] _mul_rshift_round_clip_17_rshift_source_count;
  reg [5-1:0] _mul_rshift_round_clip_17_rshift_source_mode;
  reg [16-1:0] _mul_rshift_round_clip_17_rshift_source_generator_id;
  reg [32-1:0] _mul_rshift_round_clip_17_rshift_source_offset;
  reg [33-1:0] _mul_rshift_round_clip_17_rshift_source_size;
  reg [32-1:0] _mul_rshift_round_clip_17_rshift_source_stride;
  reg [32-1:0] _mul_rshift_round_clip_17_rshift_source_offset_buf;
  reg [33-1:0] _mul_rshift_round_clip_17_rshift_source_size_buf;
  reg [32-1:0] _mul_rshift_round_clip_17_rshift_source_stride_buf;
  reg [8-1:0] _mul_rshift_round_clip_17_rshift_source_sel;
  reg [32-1:0] _mul_rshift_round_clip_17_rshift_source_ram_raddr;
  reg _mul_rshift_round_clip_17_rshift_source_ram_renable;
  wire [32-1:0] _mul_rshift_round_clip_17_rshift_source_ram_rdata;
  reg _mul_rshift_round_clip_17_rshift_source_fifo_deq;
  wire [32-1:0] _mul_rshift_round_clip_17_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_rshift_round_clip_17_rshift_source_empty_data;
  reg [33-1:0] _mul_rshift_round_clip_17_z_sink_count;
  reg [5-1:0] _mul_rshift_round_clip_17_z_sink_mode;
  reg [16-1:0] _mul_rshift_round_clip_17_z_sink_generator_id;
  reg [32-1:0] _mul_rshift_round_clip_17_z_sink_offset;
  reg [33-1:0] _mul_rshift_round_clip_17_z_sink_size;
  reg [32-1:0] _mul_rshift_round_clip_17_z_sink_stride;
  reg [32-1:0] _mul_rshift_round_clip_17_z_sink_offset_buf;
  reg [33-1:0] _mul_rshift_round_clip_17_z_sink_size_buf;
  reg [32-1:0] _mul_rshift_round_clip_17_z_sink_stride_buf;
  reg [8-1:0] _mul_rshift_round_clip_17_z_sink_sel;
  reg [32-1:0] _mul_rshift_round_clip_17_z_sink_waddr;
  reg _mul_rshift_round_clip_17_z_sink_wenable;
  reg [16-1:0] _mul_rshift_round_clip_17_z_sink_wdata;
  reg _mul_rshift_round_clip_17_z_sink_fifo_enq;
  reg [16-1:0] _mul_rshift_round_clip_17_z_sink_fifo_wdata;
  reg [16-1:0] _mul_rshift_round_clip_17_z_sink_immediate;
  reg _mul_18_stream_ivalid;
  wire _mul_18_stream_oready;
  wire _mul_18_stream_internal_oready;
  assign _mul_18_stream_internal_oready = 1;
  reg [32-1:0] _mul_18_fsm;
  localparam _mul_18_fsm_init = 0;
  wire _mul_18_run_flag;
  assign _mul_18_run_flag = 0;
  reg _mul_18_source_start;
  wire _mul_18_source_stop;
  reg _mul_18_source_busy;
  wire _mul_18_sink_start;
  wire _mul_18_sink_stop;
  wire _mul_18_sink_busy;
  wire _mul_18_busy;
  reg _mul_18_busy_reg;
  wire _mul_18_is_root;
  reg _mul_18_x_idle;
  reg [33-1:0] _mul_18_x_source_count;
  reg [5-1:0] _mul_18_x_source_mode;
  reg [16-1:0] _mul_18_x_source_generator_id;
  reg [32-1:0] _mul_18_x_source_offset;
  reg [33-1:0] _mul_18_x_source_size;
  reg [32-1:0] _mul_18_x_source_stride;
  reg [32-1:0] _mul_18_x_source_offset_buf;
  reg [33-1:0] _mul_18_x_source_size_buf;
  reg [32-1:0] _mul_18_x_source_stride_buf;
  reg [8-1:0] _mul_18_x_source_sel;
  reg [32-1:0] _mul_18_x_source_ram_raddr;
  reg _mul_18_x_source_ram_renable;
  wire [16-1:0] _mul_18_x_source_ram_rdata;
  reg _mul_18_x_source_fifo_deq;
  wire [16-1:0] _mul_18_x_source_fifo_rdata;
  reg [16-1:0] _mul_18_x_source_empty_data;
  reg _mul_18_y_idle;
  reg [33-1:0] _mul_18_y_source_count;
  reg [5-1:0] _mul_18_y_source_mode;
  reg [16-1:0] _mul_18_y_source_generator_id;
  reg [32-1:0] _mul_18_y_source_offset;
  reg [33-1:0] _mul_18_y_source_size;
  reg [32-1:0] _mul_18_y_source_stride;
  reg [32-1:0] _mul_18_y_source_offset_buf;
  reg [33-1:0] _mul_18_y_source_size_buf;
  reg [32-1:0] _mul_18_y_source_stride_buf;
  reg [8-1:0] _mul_18_y_source_sel;
  reg [32-1:0] _mul_18_y_source_ram_raddr;
  reg _mul_18_y_source_ram_renable;
  wire [16-1:0] _mul_18_y_source_ram_rdata;
  reg _mul_18_y_source_fifo_deq;
  wire [16-1:0] _mul_18_y_source_fifo_rdata;
  reg [16-1:0] _mul_18_y_source_empty_data;
  reg _mul_18_rshift_idle;
  reg [33-1:0] _mul_18_rshift_source_count;
  reg [5-1:0] _mul_18_rshift_source_mode;
  reg [16-1:0] _mul_18_rshift_source_generator_id;
  reg [32-1:0] _mul_18_rshift_source_offset;
  reg [33-1:0] _mul_18_rshift_source_size;
  reg [32-1:0] _mul_18_rshift_source_stride;
  reg [32-1:0] _mul_18_rshift_source_offset_buf;
  reg [33-1:0] _mul_18_rshift_source_size_buf;
  reg [32-1:0] _mul_18_rshift_source_stride_buf;
  reg [8-1:0] _mul_18_rshift_source_sel;
  reg [32-1:0] _mul_18_rshift_source_ram_raddr;
  reg _mul_18_rshift_source_ram_renable;
  wire [32-1:0] _mul_18_rshift_source_ram_rdata;
  reg _mul_18_rshift_source_fifo_deq;
  wire [32-1:0] _mul_18_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_18_rshift_source_empty_data;
  reg [33-1:0] _mul_18_z_sink_count;
  reg [5-1:0] _mul_18_z_sink_mode;
  reg [16-1:0] _mul_18_z_sink_generator_id;
  reg [32-1:0] _mul_18_z_sink_offset;
  reg [33-1:0] _mul_18_z_sink_size;
  reg [32-1:0] _mul_18_z_sink_stride;
  reg [32-1:0] _mul_18_z_sink_offset_buf;
  reg [33-1:0] _mul_18_z_sink_size_buf;
  reg [32-1:0] _mul_18_z_sink_stride_buf;
  reg [8-1:0] _mul_18_z_sink_sel;
  reg [32-1:0] _mul_18_z_sink_waddr;
  reg _mul_18_z_sink_wenable;
  reg [32-1:0] _mul_18_z_sink_wdata;
  reg _mul_18_z_sink_fifo_enq;
  reg [32-1:0] _mul_18_z_sink_fifo_wdata;
  reg [32-1:0] _mul_18_z_sink_immediate;
  reg _mul_19_stream_ivalid;
  wire _mul_19_stream_oready;
  wire _mul_19_stream_internal_oready;
  assign _mul_19_stream_internal_oready = 1;
  reg [32-1:0] _mul_19_fsm;
  localparam _mul_19_fsm_init = 0;
  wire _mul_19_run_flag;
  assign _mul_19_run_flag = 0;
  reg _mul_19_source_start;
  wire _mul_19_source_stop;
  reg _mul_19_source_busy;
  wire _mul_19_sink_start;
  wire _mul_19_sink_stop;
  wire _mul_19_sink_busy;
  wire _mul_19_busy;
  reg _mul_19_busy_reg;
  wire _mul_19_is_root;
  reg _mul_19_x_idle;
  reg [33-1:0] _mul_19_x_source_count;
  reg [5-1:0] _mul_19_x_source_mode;
  reg [16-1:0] _mul_19_x_source_generator_id;
  reg [32-1:0] _mul_19_x_source_offset;
  reg [33-1:0] _mul_19_x_source_size;
  reg [32-1:0] _mul_19_x_source_stride;
  reg [32-1:0] _mul_19_x_source_offset_buf;
  reg [33-1:0] _mul_19_x_source_size_buf;
  reg [32-1:0] _mul_19_x_source_stride_buf;
  reg [8-1:0] _mul_19_x_source_sel;
  reg [32-1:0] _mul_19_x_source_ram_raddr;
  reg _mul_19_x_source_ram_renable;
  wire [16-1:0] _mul_19_x_source_ram_rdata;
  reg _mul_19_x_source_fifo_deq;
  wire [16-1:0] _mul_19_x_source_fifo_rdata;
  reg [16-1:0] _mul_19_x_source_empty_data;
  reg _mul_19_y_idle;
  reg [33-1:0] _mul_19_y_source_count;
  reg [5-1:0] _mul_19_y_source_mode;
  reg [16-1:0] _mul_19_y_source_generator_id;
  reg [32-1:0] _mul_19_y_source_offset;
  reg [33-1:0] _mul_19_y_source_size;
  reg [32-1:0] _mul_19_y_source_stride;
  reg [32-1:0] _mul_19_y_source_offset_buf;
  reg [33-1:0] _mul_19_y_source_size_buf;
  reg [32-1:0] _mul_19_y_source_stride_buf;
  reg [8-1:0] _mul_19_y_source_sel;
  reg [32-1:0] _mul_19_y_source_ram_raddr;
  reg _mul_19_y_source_ram_renable;
  wire [16-1:0] _mul_19_y_source_ram_rdata;
  reg _mul_19_y_source_fifo_deq;
  wire [16-1:0] _mul_19_y_source_fifo_rdata;
  reg [16-1:0] _mul_19_y_source_empty_data;
  reg _mul_19_rshift_idle;
  reg [33-1:0] _mul_19_rshift_source_count;
  reg [5-1:0] _mul_19_rshift_source_mode;
  reg [16-1:0] _mul_19_rshift_source_generator_id;
  reg [32-1:0] _mul_19_rshift_source_offset;
  reg [33-1:0] _mul_19_rshift_source_size;
  reg [32-1:0] _mul_19_rshift_source_stride;
  reg [32-1:0] _mul_19_rshift_source_offset_buf;
  reg [33-1:0] _mul_19_rshift_source_size_buf;
  reg [32-1:0] _mul_19_rshift_source_stride_buf;
  reg [8-1:0] _mul_19_rshift_source_sel;
  reg [32-1:0] _mul_19_rshift_source_ram_raddr;
  reg _mul_19_rshift_source_ram_renable;
  wire [32-1:0] _mul_19_rshift_source_ram_rdata;
  reg _mul_19_rshift_source_fifo_deq;
  wire [32-1:0] _mul_19_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_19_rshift_source_empty_data;
  reg [33-1:0] _mul_19_z_sink_count;
  reg [5-1:0] _mul_19_z_sink_mode;
  reg [16-1:0] _mul_19_z_sink_generator_id;
  reg [32-1:0] _mul_19_z_sink_offset;
  reg [33-1:0] _mul_19_z_sink_size;
  reg [32-1:0] _mul_19_z_sink_stride;
  reg [32-1:0] _mul_19_z_sink_offset_buf;
  reg [33-1:0] _mul_19_z_sink_size_buf;
  reg [32-1:0] _mul_19_z_sink_stride_buf;
  reg [8-1:0] _mul_19_z_sink_sel;
  reg [32-1:0] _mul_19_z_sink_waddr;
  reg _mul_19_z_sink_wenable;
  reg [32-1:0] _mul_19_z_sink_wdata;
  reg _mul_19_z_sink_fifo_enq;
  reg [32-1:0] _mul_19_z_sink_fifo_wdata;
  reg [32-1:0] _mul_19_z_sink_immediate;
  reg _mul_20_stream_ivalid;
  wire _mul_20_stream_oready;
  wire _mul_20_stream_internal_oready;
  assign _mul_20_stream_internal_oready = 1;
  reg [32-1:0] _mul_20_fsm;
  localparam _mul_20_fsm_init = 0;
  wire _mul_20_run_flag;
  assign _mul_20_run_flag = 0;
  reg _mul_20_source_start;
  wire _mul_20_source_stop;
  reg _mul_20_source_busy;
  wire _mul_20_sink_start;
  wire _mul_20_sink_stop;
  wire _mul_20_sink_busy;
  wire _mul_20_busy;
  reg _mul_20_busy_reg;
  wire _mul_20_is_root;
  reg _mul_20_x_idle;
  reg [33-1:0] _mul_20_x_source_count;
  reg [5-1:0] _mul_20_x_source_mode;
  reg [16-1:0] _mul_20_x_source_generator_id;
  reg [32-1:0] _mul_20_x_source_offset;
  reg [33-1:0] _mul_20_x_source_size;
  reg [32-1:0] _mul_20_x_source_stride;
  reg [32-1:0] _mul_20_x_source_offset_buf;
  reg [33-1:0] _mul_20_x_source_size_buf;
  reg [32-1:0] _mul_20_x_source_stride_buf;
  reg [8-1:0] _mul_20_x_source_sel;
  reg [32-1:0] _mul_20_x_source_ram_raddr;
  reg _mul_20_x_source_ram_renable;
  wire [16-1:0] _mul_20_x_source_ram_rdata;
  reg _mul_20_x_source_fifo_deq;
  wire [16-1:0] _mul_20_x_source_fifo_rdata;
  reg [16-1:0] _mul_20_x_source_empty_data;
  reg _mul_20_y_idle;
  reg [33-1:0] _mul_20_y_source_count;
  reg [5-1:0] _mul_20_y_source_mode;
  reg [16-1:0] _mul_20_y_source_generator_id;
  reg [32-1:0] _mul_20_y_source_offset;
  reg [33-1:0] _mul_20_y_source_size;
  reg [32-1:0] _mul_20_y_source_stride;
  reg [32-1:0] _mul_20_y_source_offset_buf;
  reg [33-1:0] _mul_20_y_source_size_buf;
  reg [32-1:0] _mul_20_y_source_stride_buf;
  reg [8-1:0] _mul_20_y_source_sel;
  reg [32-1:0] _mul_20_y_source_ram_raddr;
  reg _mul_20_y_source_ram_renable;
  wire [16-1:0] _mul_20_y_source_ram_rdata;
  reg _mul_20_y_source_fifo_deq;
  wire [16-1:0] _mul_20_y_source_fifo_rdata;
  reg [16-1:0] _mul_20_y_source_empty_data;
  reg _mul_20_rshift_idle;
  reg [33-1:0] _mul_20_rshift_source_count;
  reg [5-1:0] _mul_20_rshift_source_mode;
  reg [16-1:0] _mul_20_rshift_source_generator_id;
  reg [32-1:0] _mul_20_rshift_source_offset;
  reg [33-1:0] _mul_20_rshift_source_size;
  reg [32-1:0] _mul_20_rshift_source_stride;
  reg [32-1:0] _mul_20_rshift_source_offset_buf;
  reg [33-1:0] _mul_20_rshift_source_size_buf;
  reg [32-1:0] _mul_20_rshift_source_stride_buf;
  reg [8-1:0] _mul_20_rshift_source_sel;
  reg [32-1:0] _mul_20_rshift_source_ram_raddr;
  reg _mul_20_rshift_source_ram_renable;
  wire [32-1:0] _mul_20_rshift_source_ram_rdata;
  reg _mul_20_rshift_source_fifo_deq;
  wire [32-1:0] _mul_20_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_20_rshift_source_empty_data;
  reg [33-1:0] _mul_20_z_sink_count;
  reg [5-1:0] _mul_20_z_sink_mode;
  reg [16-1:0] _mul_20_z_sink_generator_id;
  reg [32-1:0] _mul_20_z_sink_offset;
  reg [33-1:0] _mul_20_z_sink_size;
  reg [32-1:0] _mul_20_z_sink_stride;
  reg [32-1:0] _mul_20_z_sink_offset_buf;
  reg [33-1:0] _mul_20_z_sink_size_buf;
  reg [32-1:0] _mul_20_z_sink_stride_buf;
  reg [8-1:0] _mul_20_z_sink_sel;
  reg [32-1:0] _mul_20_z_sink_waddr;
  reg _mul_20_z_sink_wenable;
  reg [32-1:0] _mul_20_z_sink_wdata;
  reg _mul_20_z_sink_fifo_enq;
  reg [32-1:0] _mul_20_z_sink_fifo_wdata;
  reg [32-1:0] _mul_20_z_sink_immediate;
  reg _mul_21_stream_ivalid;
  wire _mul_21_stream_oready;
  wire _mul_21_stream_internal_oready;
  assign _mul_21_stream_internal_oready = 1;
  reg [32-1:0] _mul_21_fsm;
  localparam _mul_21_fsm_init = 0;
  wire _mul_21_run_flag;
  assign _mul_21_run_flag = 0;
  reg _mul_21_source_start;
  wire _mul_21_source_stop;
  reg _mul_21_source_busy;
  wire _mul_21_sink_start;
  wire _mul_21_sink_stop;
  wire _mul_21_sink_busy;
  wire _mul_21_busy;
  reg _mul_21_busy_reg;
  wire _mul_21_is_root;
  reg _mul_21_x_idle;
  reg [33-1:0] _mul_21_x_source_count;
  reg [5-1:0] _mul_21_x_source_mode;
  reg [16-1:0] _mul_21_x_source_generator_id;
  reg [32-1:0] _mul_21_x_source_offset;
  reg [33-1:0] _mul_21_x_source_size;
  reg [32-1:0] _mul_21_x_source_stride;
  reg [32-1:0] _mul_21_x_source_offset_buf;
  reg [33-1:0] _mul_21_x_source_size_buf;
  reg [32-1:0] _mul_21_x_source_stride_buf;
  reg [8-1:0] _mul_21_x_source_sel;
  reg [32-1:0] _mul_21_x_source_ram_raddr;
  reg _mul_21_x_source_ram_renable;
  wire [16-1:0] _mul_21_x_source_ram_rdata;
  reg _mul_21_x_source_fifo_deq;
  wire [16-1:0] _mul_21_x_source_fifo_rdata;
  reg [16-1:0] _mul_21_x_source_empty_data;
  reg _mul_21_y_idle;
  reg [33-1:0] _mul_21_y_source_count;
  reg [5-1:0] _mul_21_y_source_mode;
  reg [16-1:0] _mul_21_y_source_generator_id;
  reg [32-1:0] _mul_21_y_source_offset;
  reg [33-1:0] _mul_21_y_source_size;
  reg [32-1:0] _mul_21_y_source_stride;
  reg [32-1:0] _mul_21_y_source_offset_buf;
  reg [33-1:0] _mul_21_y_source_size_buf;
  reg [32-1:0] _mul_21_y_source_stride_buf;
  reg [8-1:0] _mul_21_y_source_sel;
  reg [32-1:0] _mul_21_y_source_ram_raddr;
  reg _mul_21_y_source_ram_renable;
  wire [16-1:0] _mul_21_y_source_ram_rdata;
  reg _mul_21_y_source_fifo_deq;
  wire [16-1:0] _mul_21_y_source_fifo_rdata;
  reg [16-1:0] _mul_21_y_source_empty_data;
  reg _mul_21_rshift_idle;
  reg [33-1:0] _mul_21_rshift_source_count;
  reg [5-1:0] _mul_21_rshift_source_mode;
  reg [16-1:0] _mul_21_rshift_source_generator_id;
  reg [32-1:0] _mul_21_rshift_source_offset;
  reg [33-1:0] _mul_21_rshift_source_size;
  reg [32-1:0] _mul_21_rshift_source_stride;
  reg [32-1:0] _mul_21_rshift_source_offset_buf;
  reg [33-1:0] _mul_21_rshift_source_size_buf;
  reg [32-1:0] _mul_21_rshift_source_stride_buf;
  reg [8-1:0] _mul_21_rshift_source_sel;
  reg [32-1:0] _mul_21_rshift_source_ram_raddr;
  reg _mul_21_rshift_source_ram_renable;
  wire [32-1:0] _mul_21_rshift_source_ram_rdata;
  reg _mul_21_rshift_source_fifo_deq;
  wire [32-1:0] _mul_21_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_21_rshift_source_empty_data;
  reg [33-1:0] _mul_21_z_sink_count;
  reg [5-1:0] _mul_21_z_sink_mode;
  reg [16-1:0] _mul_21_z_sink_generator_id;
  reg [32-1:0] _mul_21_z_sink_offset;
  reg [33-1:0] _mul_21_z_sink_size;
  reg [32-1:0] _mul_21_z_sink_stride;
  reg [32-1:0] _mul_21_z_sink_offset_buf;
  reg [33-1:0] _mul_21_z_sink_size_buf;
  reg [32-1:0] _mul_21_z_sink_stride_buf;
  reg [8-1:0] _mul_21_z_sink_sel;
  reg [32-1:0] _mul_21_z_sink_waddr;
  reg _mul_21_z_sink_wenable;
  reg [32-1:0] _mul_21_z_sink_wdata;
  reg _mul_21_z_sink_fifo_enq;
  reg [32-1:0] _mul_21_z_sink_fifo_wdata;
  reg [32-1:0] _mul_21_z_sink_immediate;
  reg _mul_22_stream_ivalid;
  wire _mul_22_stream_oready;
  wire _mul_22_stream_internal_oready;
  assign _mul_22_stream_internal_oready = 1;
  reg [32-1:0] _mul_22_fsm;
  localparam _mul_22_fsm_init = 0;
  wire _mul_22_run_flag;
  assign _mul_22_run_flag = 0;
  reg _mul_22_source_start;
  wire _mul_22_source_stop;
  reg _mul_22_source_busy;
  wire _mul_22_sink_start;
  wire _mul_22_sink_stop;
  wire _mul_22_sink_busy;
  wire _mul_22_busy;
  reg _mul_22_busy_reg;
  wire _mul_22_is_root;
  reg _mul_22_x_idle;
  reg [33-1:0] _mul_22_x_source_count;
  reg [5-1:0] _mul_22_x_source_mode;
  reg [16-1:0] _mul_22_x_source_generator_id;
  reg [32-1:0] _mul_22_x_source_offset;
  reg [33-1:0] _mul_22_x_source_size;
  reg [32-1:0] _mul_22_x_source_stride;
  reg [32-1:0] _mul_22_x_source_offset_buf;
  reg [33-1:0] _mul_22_x_source_size_buf;
  reg [32-1:0] _mul_22_x_source_stride_buf;
  reg [8-1:0] _mul_22_x_source_sel;
  reg [32-1:0] _mul_22_x_source_ram_raddr;
  reg _mul_22_x_source_ram_renable;
  wire [16-1:0] _mul_22_x_source_ram_rdata;
  reg _mul_22_x_source_fifo_deq;
  wire [16-1:0] _mul_22_x_source_fifo_rdata;
  reg [16-1:0] _mul_22_x_source_empty_data;
  reg _mul_22_y_idle;
  reg [33-1:0] _mul_22_y_source_count;
  reg [5-1:0] _mul_22_y_source_mode;
  reg [16-1:0] _mul_22_y_source_generator_id;
  reg [32-1:0] _mul_22_y_source_offset;
  reg [33-1:0] _mul_22_y_source_size;
  reg [32-1:0] _mul_22_y_source_stride;
  reg [32-1:0] _mul_22_y_source_offset_buf;
  reg [33-1:0] _mul_22_y_source_size_buf;
  reg [32-1:0] _mul_22_y_source_stride_buf;
  reg [8-1:0] _mul_22_y_source_sel;
  reg [32-1:0] _mul_22_y_source_ram_raddr;
  reg _mul_22_y_source_ram_renable;
  wire [16-1:0] _mul_22_y_source_ram_rdata;
  reg _mul_22_y_source_fifo_deq;
  wire [16-1:0] _mul_22_y_source_fifo_rdata;
  reg [16-1:0] _mul_22_y_source_empty_data;
  reg _mul_22_rshift_idle;
  reg [33-1:0] _mul_22_rshift_source_count;
  reg [5-1:0] _mul_22_rshift_source_mode;
  reg [16-1:0] _mul_22_rshift_source_generator_id;
  reg [32-1:0] _mul_22_rshift_source_offset;
  reg [33-1:0] _mul_22_rshift_source_size;
  reg [32-1:0] _mul_22_rshift_source_stride;
  reg [32-1:0] _mul_22_rshift_source_offset_buf;
  reg [33-1:0] _mul_22_rshift_source_size_buf;
  reg [32-1:0] _mul_22_rshift_source_stride_buf;
  reg [8-1:0] _mul_22_rshift_source_sel;
  reg [32-1:0] _mul_22_rshift_source_ram_raddr;
  reg _mul_22_rshift_source_ram_renable;
  wire [32-1:0] _mul_22_rshift_source_ram_rdata;
  reg _mul_22_rshift_source_fifo_deq;
  wire [32-1:0] _mul_22_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_22_rshift_source_empty_data;
  reg [33-1:0] _mul_22_z_sink_count;
  reg [5-1:0] _mul_22_z_sink_mode;
  reg [16-1:0] _mul_22_z_sink_generator_id;
  reg [32-1:0] _mul_22_z_sink_offset;
  reg [33-1:0] _mul_22_z_sink_size;
  reg [32-1:0] _mul_22_z_sink_stride;
  reg [32-1:0] _mul_22_z_sink_offset_buf;
  reg [33-1:0] _mul_22_z_sink_size_buf;
  reg [32-1:0] _mul_22_z_sink_stride_buf;
  reg [8-1:0] _mul_22_z_sink_sel;
  reg [32-1:0] _mul_22_z_sink_waddr;
  reg _mul_22_z_sink_wenable;
  reg [32-1:0] _mul_22_z_sink_wdata;
  reg _mul_22_z_sink_fifo_enq;
  reg [32-1:0] _mul_22_z_sink_fifo_wdata;
  reg [32-1:0] _mul_22_z_sink_immediate;
  reg _mul_23_stream_ivalid;
  wire _mul_23_stream_oready;
  wire _mul_23_stream_internal_oready;
  assign _mul_23_stream_internal_oready = 1;
  reg [32-1:0] _mul_23_fsm;
  localparam _mul_23_fsm_init = 0;
  wire _mul_23_run_flag;
  assign _mul_23_run_flag = 0;
  reg _mul_23_source_start;
  wire _mul_23_source_stop;
  reg _mul_23_source_busy;
  wire _mul_23_sink_start;
  wire _mul_23_sink_stop;
  wire _mul_23_sink_busy;
  wire _mul_23_busy;
  reg _mul_23_busy_reg;
  wire _mul_23_is_root;
  reg _mul_23_x_idle;
  reg [33-1:0] _mul_23_x_source_count;
  reg [5-1:0] _mul_23_x_source_mode;
  reg [16-1:0] _mul_23_x_source_generator_id;
  reg [32-1:0] _mul_23_x_source_offset;
  reg [33-1:0] _mul_23_x_source_size;
  reg [32-1:0] _mul_23_x_source_stride;
  reg [32-1:0] _mul_23_x_source_offset_buf;
  reg [33-1:0] _mul_23_x_source_size_buf;
  reg [32-1:0] _mul_23_x_source_stride_buf;
  reg [8-1:0] _mul_23_x_source_sel;
  reg [32-1:0] _mul_23_x_source_ram_raddr;
  reg _mul_23_x_source_ram_renable;
  wire [16-1:0] _mul_23_x_source_ram_rdata;
  reg _mul_23_x_source_fifo_deq;
  wire [16-1:0] _mul_23_x_source_fifo_rdata;
  reg [16-1:0] _mul_23_x_source_empty_data;
  reg _mul_23_y_idle;
  reg [33-1:0] _mul_23_y_source_count;
  reg [5-1:0] _mul_23_y_source_mode;
  reg [16-1:0] _mul_23_y_source_generator_id;
  reg [32-1:0] _mul_23_y_source_offset;
  reg [33-1:0] _mul_23_y_source_size;
  reg [32-1:0] _mul_23_y_source_stride;
  reg [32-1:0] _mul_23_y_source_offset_buf;
  reg [33-1:0] _mul_23_y_source_size_buf;
  reg [32-1:0] _mul_23_y_source_stride_buf;
  reg [8-1:0] _mul_23_y_source_sel;
  reg [32-1:0] _mul_23_y_source_ram_raddr;
  reg _mul_23_y_source_ram_renable;
  wire [16-1:0] _mul_23_y_source_ram_rdata;
  reg _mul_23_y_source_fifo_deq;
  wire [16-1:0] _mul_23_y_source_fifo_rdata;
  reg [16-1:0] _mul_23_y_source_empty_data;
  reg _mul_23_rshift_idle;
  reg [33-1:0] _mul_23_rshift_source_count;
  reg [5-1:0] _mul_23_rshift_source_mode;
  reg [16-1:0] _mul_23_rshift_source_generator_id;
  reg [32-1:0] _mul_23_rshift_source_offset;
  reg [33-1:0] _mul_23_rshift_source_size;
  reg [32-1:0] _mul_23_rshift_source_stride;
  reg [32-1:0] _mul_23_rshift_source_offset_buf;
  reg [33-1:0] _mul_23_rshift_source_size_buf;
  reg [32-1:0] _mul_23_rshift_source_stride_buf;
  reg [8-1:0] _mul_23_rshift_source_sel;
  reg [32-1:0] _mul_23_rshift_source_ram_raddr;
  reg _mul_23_rshift_source_ram_renable;
  wire [32-1:0] _mul_23_rshift_source_ram_rdata;
  reg _mul_23_rshift_source_fifo_deq;
  wire [32-1:0] _mul_23_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_23_rshift_source_empty_data;
  reg [33-1:0] _mul_23_z_sink_count;
  reg [5-1:0] _mul_23_z_sink_mode;
  reg [16-1:0] _mul_23_z_sink_generator_id;
  reg [32-1:0] _mul_23_z_sink_offset;
  reg [33-1:0] _mul_23_z_sink_size;
  reg [32-1:0] _mul_23_z_sink_stride;
  reg [32-1:0] _mul_23_z_sink_offset_buf;
  reg [33-1:0] _mul_23_z_sink_size_buf;
  reg [32-1:0] _mul_23_z_sink_stride_buf;
  reg [8-1:0] _mul_23_z_sink_sel;
  reg [32-1:0] _mul_23_z_sink_waddr;
  reg _mul_23_z_sink_wenable;
  reg [32-1:0] _mul_23_z_sink_wdata;
  reg _mul_23_z_sink_fifo_enq;
  reg [32-1:0] _mul_23_z_sink_fifo_wdata;
  reg [32-1:0] _mul_23_z_sink_immediate;
  reg _mul_24_stream_ivalid;
  wire _mul_24_stream_oready;
  wire _mul_24_stream_internal_oready;
  assign _mul_24_stream_internal_oready = 1;
  reg [32-1:0] _mul_24_fsm;
  localparam _mul_24_fsm_init = 0;
  wire _mul_24_run_flag;
  assign _mul_24_run_flag = 0;
  reg _mul_24_source_start;
  wire _mul_24_source_stop;
  reg _mul_24_source_busy;
  wire _mul_24_sink_start;
  wire _mul_24_sink_stop;
  wire _mul_24_sink_busy;
  wire _mul_24_busy;
  reg _mul_24_busy_reg;
  wire _mul_24_is_root;
  reg _mul_24_x_idle;
  reg [33-1:0] _mul_24_x_source_count;
  reg [5-1:0] _mul_24_x_source_mode;
  reg [16-1:0] _mul_24_x_source_generator_id;
  reg [32-1:0] _mul_24_x_source_offset;
  reg [33-1:0] _mul_24_x_source_size;
  reg [32-1:0] _mul_24_x_source_stride;
  reg [32-1:0] _mul_24_x_source_offset_buf;
  reg [33-1:0] _mul_24_x_source_size_buf;
  reg [32-1:0] _mul_24_x_source_stride_buf;
  reg [8-1:0] _mul_24_x_source_sel;
  reg [32-1:0] _mul_24_x_source_ram_raddr;
  reg _mul_24_x_source_ram_renable;
  wire [16-1:0] _mul_24_x_source_ram_rdata;
  reg _mul_24_x_source_fifo_deq;
  wire [16-1:0] _mul_24_x_source_fifo_rdata;
  reg [16-1:0] _mul_24_x_source_empty_data;
  reg _mul_24_y_idle;
  reg [33-1:0] _mul_24_y_source_count;
  reg [5-1:0] _mul_24_y_source_mode;
  reg [16-1:0] _mul_24_y_source_generator_id;
  reg [32-1:0] _mul_24_y_source_offset;
  reg [33-1:0] _mul_24_y_source_size;
  reg [32-1:0] _mul_24_y_source_stride;
  reg [32-1:0] _mul_24_y_source_offset_buf;
  reg [33-1:0] _mul_24_y_source_size_buf;
  reg [32-1:0] _mul_24_y_source_stride_buf;
  reg [8-1:0] _mul_24_y_source_sel;
  reg [32-1:0] _mul_24_y_source_ram_raddr;
  reg _mul_24_y_source_ram_renable;
  wire [16-1:0] _mul_24_y_source_ram_rdata;
  reg _mul_24_y_source_fifo_deq;
  wire [16-1:0] _mul_24_y_source_fifo_rdata;
  reg [16-1:0] _mul_24_y_source_empty_data;
  reg _mul_24_rshift_idle;
  reg [33-1:0] _mul_24_rshift_source_count;
  reg [5-1:0] _mul_24_rshift_source_mode;
  reg [16-1:0] _mul_24_rshift_source_generator_id;
  reg [32-1:0] _mul_24_rshift_source_offset;
  reg [33-1:0] _mul_24_rshift_source_size;
  reg [32-1:0] _mul_24_rshift_source_stride;
  reg [32-1:0] _mul_24_rshift_source_offset_buf;
  reg [33-1:0] _mul_24_rshift_source_size_buf;
  reg [32-1:0] _mul_24_rshift_source_stride_buf;
  reg [8-1:0] _mul_24_rshift_source_sel;
  reg [32-1:0] _mul_24_rshift_source_ram_raddr;
  reg _mul_24_rshift_source_ram_renable;
  wire [32-1:0] _mul_24_rshift_source_ram_rdata;
  reg _mul_24_rshift_source_fifo_deq;
  wire [32-1:0] _mul_24_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_24_rshift_source_empty_data;
  reg [33-1:0] _mul_24_z_sink_count;
  reg [5-1:0] _mul_24_z_sink_mode;
  reg [16-1:0] _mul_24_z_sink_generator_id;
  reg [32-1:0] _mul_24_z_sink_offset;
  reg [33-1:0] _mul_24_z_sink_size;
  reg [32-1:0] _mul_24_z_sink_stride;
  reg [32-1:0] _mul_24_z_sink_offset_buf;
  reg [33-1:0] _mul_24_z_sink_size_buf;
  reg [32-1:0] _mul_24_z_sink_stride_buf;
  reg [8-1:0] _mul_24_z_sink_sel;
  reg [32-1:0] _mul_24_z_sink_waddr;
  reg _mul_24_z_sink_wenable;
  reg [32-1:0] _mul_24_z_sink_wdata;
  reg _mul_24_z_sink_fifo_enq;
  reg [32-1:0] _mul_24_z_sink_fifo_wdata;
  reg [32-1:0] _mul_24_z_sink_immediate;
  reg _mul_25_stream_ivalid;
  wire _mul_25_stream_oready;
  wire _mul_25_stream_internal_oready;
  assign _mul_25_stream_internal_oready = 1;
  reg [32-1:0] _mul_25_fsm;
  localparam _mul_25_fsm_init = 0;
  wire _mul_25_run_flag;
  assign _mul_25_run_flag = 0;
  reg _mul_25_source_start;
  wire _mul_25_source_stop;
  reg _mul_25_source_busy;
  wire _mul_25_sink_start;
  wire _mul_25_sink_stop;
  wire _mul_25_sink_busy;
  wire _mul_25_busy;
  reg _mul_25_busy_reg;
  wire _mul_25_is_root;
  reg _mul_25_x_idle;
  reg [33-1:0] _mul_25_x_source_count;
  reg [5-1:0] _mul_25_x_source_mode;
  reg [16-1:0] _mul_25_x_source_generator_id;
  reg [32-1:0] _mul_25_x_source_offset;
  reg [33-1:0] _mul_25_x_source_size;
  reg [32-1:0] _mul_25_x_source_stride;
  reg [32-1:0] _mul_25_x_source_offset_buf;
  reg [33-1:0] _mul_25_x_source_size_buf;
  reg [32-1:0] _mul_25_x_source_stride_buf;
  reg [8-1:0] _mul_25_x_source_sel;
  reg [32-1:0] _mul_25_x_source_ram_raddr;
  reg _mul_25_x_source_ram_renable;
  wire [16-1:0] _mul_25_x_source_ram_rdata;
  reg _mul_25_x_source_fifo_deq;
  wire [16-1:0] _mul_25_x_source_fifo_rdata;
  reg [16-1:0] _mul_25_x_source_empty_data;
  reg _mul_25_y_idle;
  reg [33-1:0] _mul_25_y_source_count;
  reg [5-1:0] _mul_25_y_source_mode;
  reg [16-1:0] _mul_25_y_source_generator_id;
  reg [32-1:0] _mul_25_y_source_offset;
  reg [33-1:0] _mul_25_y_source_size;
  reg [32-1:0] _mul_25_y_source_stride;
  reg [32-1:0] _mul_25_y_source_offset_buf;
  reg [33-1:0] _mul_25_y_source_size_buf;
  reg [32-1:0] _mul_25_y_source_stride_buf;
  reg [8-1:0] _mul_25_y_source_sel;
  reg [32-1:0] _mul_25_y_source_ram_raddr;
  reg _mul_25_y_source_ram_renable;
  wire [16-1:0] _mul_25_y_source_ram_rdata;
  reg _mul_25_y_source_fifo_deq;
  wire [16-1:0] _mul_25_y_source_fifo_rdata;
  reg [16-1:0] _mul_25_y_source_empty_data;
  reg _mul_25_rshift_idle;
  reg [33-1:0] _mul_25_rshift_source_count;
  reg [5-1:0] _mul_25_rshift_source_mode;
  reg [16-1:0] _mul_25_rshift_source_generator_id;
  reg [32-1:0] _mul_25_rshift_source_offset;
  reg [33-1:0] _mul_25_rshift_source_size;
  reg [32-1:0] _mul_25_rshift_source_stride;
  reg [32-1:0] _mul_25_rshift_source_offset_buf;
  reg [33-1:0] _mul_25_rshift_source_size_buf;
  reg [32-1:0] _mul_25_rshift_source_stride_buf;
  reg [8-1:0] _mul_25_rshift_source_sel;
  reg [32-1:0] _mul_25_rshift_source_ram_raddr;
  reg _mul_25_rshift_source_ram_renable;
  wire [32-1:0] _mul_25_rshift_source_ram_rdata;
  reg _mul_25_rshift_source_fifo_deq;
  wire [32-1:0] _mul_25_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_25_rshift_source_empty_data;
  reg [33-1:0] _mul_25_z_sink_count;
  reg [5-1:0] _mul_25_z_sink_mode;
  reg [16-1:0] _mul_25_z_sink_generator_id;
  reg [32-1:0] _mul_25_z_sink_offset;
  reg [33-1:0] _mul_25_z_sink_size;
  reg [32-1:0] _mul_25_z_sink_stride;
  reg [32-1:0] _mul_25_z_sink_offset_buf;
  reg [33-1:0] _mul_25_z_sink_size_buf;
  reg [32-1:0] _mul_25_z_sink_stride_buf;
  reg [8-1:0] _mul_25_z_sink_sel;
  reg [32-1:0] _mul_25_z_sink_waddr;
  reg _mul_25_z_sink_wenable;
  reg [32-1:0] _mul_25_z_sink_wdata;
  reg _mul_25_z_sink_fifo_enq;
  reg [32-1:0] _mul_25_z_sink_fifo_wdata;
  reg [32-1:0] _mul_25_z_sink_immediate;
  reg _mul_26_stream_ivalid;
  wire _mul_26_stream_oready;
  wire _mul_26_stream_internal_oready;
  assign _mul_26_stream_internal_oready = 1;
  reg [32-1:0] _mul_26_fsm;
  localparam _mul_26_fsm_init = 0;
  wire _mul_26_run_flag;
  assign _mul_26_run_flag = 0;
  reg _mul_26_source_start;
  wire _mul_26_source_stop;
  reg _mul_26_source_busy;
  wire _mul_26_sink_start;
  wire _mul_26_sink_stop;
  wire _mul_26_sink_busy;
  wire _mul_26_busy;
  reg _mul_26_busy_reg;
  wire _mul_26_is_root;
  reg _mul_26_x_idle;
  reg [33-1:0] _mul_26_x_source_count;
  reg [5-1:0] _mul_26_x_source_mode;
  reg [16-1:0] _mul_26_x_source_generator_id;
  reg [32-1:0] _mul_26_x_source_offset;
  reg [33-1:0] _mul_26_x_source_size;
  reg [32-1:0] _mul_26_x_source_stride;
  reg [32-1:0] _mul_26_x_source_offset_buf;
  reg [33-1:0] _mul_26_x_source_size_buf;
  reg [32-1:0] _mul_26_x_source_stride_buf;
  reg [8-1:0] _mul_26_x_source_sel;
  reg [32-1:0] _mul_26_x_source_ram_raddr;
  reg _mul_26_x_source_ram_renable;
  wire [16-1:0] _mul_26_x_source_ram_rdata;
  reg _mul_26_x_source_fifo_deq;
  wire [16-1:0] _mul_26_x_source_fifo_rdata;
  reg [16-1:0] _mul_26_x_source_empty_data;
  reg _mul_26_y_idle;
  reg [33-1:0] _mul_26_y_source_count;
  reg [5-1:0] _mul_26_y_source_mode;
  reg [16-1:0] _mul_26_y_source_generator_id;
  reg [32-1:0] _mul_26_y_source_offset;
  reg [33-1:0] _mul_26_y_source_size;
  reg [32-1:0] _mul_26_y_source_stride;
  reg [32-1:0] _mul_26_y_source_offset_buf;
  reg [33-1:0] _mul_26_y_source_size_buf;
  reg [32-1:0] _mul_26_y_source_stride_buf;
  reg [8-1:0] _mul_26_y_source_sel;
  reg [32-1:0] _mul_26_y_source_ram_raddr;
  reg _mul_26_y_source_ram_renable;
  wire [16-1:0] _mul_26_y_source_ram_rdata;
  reg _mul_26_y_source_fifo_deq;
  wire [16-1:0] _mul_26_y_source_fifo_rdata;
  reg [16-1:0] _mul_26_y_source_empty_data;
  reg _mul_26_rshift_idle;
  reg [33-1:0] _mul_26_rshift_source_count;
  reg [5-1:0] _mul_26_rshift_source_mode;
  reg [16-1:0] _mul_26_rshift_source_generator_id;
  reg [32-1:0] _mul_26_rshift_source_offset;
  reg [33-1:0] _mul_26_rshift_source_size;
  reg [32-1:0] _mul_26_rshift_source_stride;
  reg [32-1:0] _mul_26_rshift_source_offset_buf;
  reg [33-1:0] _mul_26_rshift_source_size_buf;
  reg [32-1:0] _mul_26_rshift_source_stride_buf;
  reg [8-1:0] _mul_26_rshift_source_sel;
  reg [32-1:0] _mul_26_rshift_source_ram_raddr;
  reg _mul_26_rshift_source_ram_renable;
  wire [32-1:0] _mul_26_rshift_source_ram_rdata;
  reg _mul_26_rshift_source_fifo_deq;
  wire [32-1:0] _mul_26_rshift_source_fifo_rdata;
  reg [32-1:0] _mul_26_rshift_source_empty_data;
  reg [33-1:0] _mul_26_z_sink_count;
  reg [5-1:0] _mul_26_z_sink_mode;
  reg [16-1:0] _mul_26_z_sink_generator_id;
  reg [32-1:0] _mul_26_z_sink_offset;
  reg [33-1:0] _mul_26_z_sink_size;
  reg [32-1:0] _mul_26_z_sink_stride;
  reg [32-1:0] _mul_26_z_sink_offset_buf;
  reg [33-1:0] _mul_26_z_sink_size_buf;
  reg [32-1:0] _mul_26_z_sink_stride_buf;
  reg [8-1:0] _mul_26_z_sink_sel;
  reg [32-1:0] _mul_26_z_sink_waddr;
  reg _mul_26_z_sink_wenable;
  reg [32-1:0] _mul_26_z_sink_wdata;
  reg _mul_26_z_sink_fifo_enq;
  reg [32-1:0] _mul_26_z_sink_fifo_wdata;
  reg [32-1:0] _mul_26_z_sink_immediate;
  reg __reduce_max_27_stream_ivalid;
  wire __reduce_max_27_stream_oready;
  wire __reduce_max_27_stream_internal_oready;
  assign __reduce_max_27_stream_internal_oready = 1;
  reg [32-1:0] __reduce_max_27_fsm;
  localparam __reduce_max_27_fsm_init = 0;
  wire __reduce_max_27_run_flag;
  assign __reduce_max_27_run_flag = 0;
  reg __reduce_max_27_source_start;
  wire __reduce_max_27_source_stop;
  reg __reduce_max_27_source_busy;
  wire __reduce_max_27_sink_start;
  wire __reduce_max_27_sink_stop;
  wire __reduce_max_27_sink_busy;
  wire __reduce_max_27_busy;
  reg __reduce_max_27_busy_reg;
  wire __reduce_max_27_is_root;
  reg __reduce_max_27_x_idle;
  reg [33-1:0] __reduce_max_27_x_source_count;
  reg [5-1:0] __reduce_max_27_x_source_mode;
  reg [16-1:0] __reduce_max_27_x_source_generator_id;
  reg [32-1:0] __reduce_max_27_x_source_offset;
  reg [33-1:0] __reduce_max_27_x_source_size;
  reg [32-1:0] __reduce_max_27_x_source_stride;
  reg [32-1:0] __reduce_max_27_x_source_offset_buf;
  reg [33-1:0] __reduce_max_27_x_source_size_buf;
  reg [32-1:0] __reduce_max_27_x_source_stride_buf;
  reg [8-1:0] __reduce_max_27_x_source_sel;
  reg [32-1:0] __reduce_max_27_x_source_ram_raddr;
  reg __reduce_max_27_x_source_ram_renable;
  wire [16-1:0] __reduce_max_27_x_source_ram_rdata;
  reg __reduce_max_27_x_source_fifo_deq;
  wire [16-1:0] __reduce_max_27_x_source_fifo_rdata;
  reg [16-1:0] __reduce_max_27_x_source_empty_data;
  reg [32-1:0] __reduce_max_27_size_next_parameter_data;
  reg [33-1:0] __reduce_max_27_data_sink_count;
  reg [5-1:0] __reduce_max_27_data_sink_mode;
  reg [16-1:0] __reduce_max_27_data_sink_generator_id;
  reg [32-1:0] __reduce_max_27_data_sink_offset;
  reg [33-1:0] __reduce_max_27_data_sink_size;
  reg [32-1:0] __reduce_max_27_data_sink_stride;
  reg [32-1:0] __reduce_max_27_data_sink_offset_buf;
  reg [33-1:0] __reduce_max_27_data_sink_size_buf;
  reg [32-1:0] __reduce_max_27_data_sink_stride_buf;
  reg [8-1:0] __reduce_max_27_data_sink_sel;
  reg [32-1:0] __reduce_max_27_data_sink_waddr;
  reg __reduce_max_27_data_sink_wenable;
  reg [16-1:0] __reduce_max_27_data_sink_wdata;
  reg __reduce_max_27_data_sink_fifo_enq;
  reg [16-1:0] __reduce_max_27_data_sink_fifo_wdata;
  reg [16-1:0] __reduce_max_27_data_sink_immediate;
  reg [33-1:0] __reduce_max_27_valid_sink_count;
  reg [5-1:0] __reduce_max_27_valid_sink_mode;
  reg [16-1:0] __reduce_max_27_valid_sink_generator_id;
  reg [32-1:0] __reduce_max_27_valid_sink_offset;
  reg [33-1:0] __reduce_max_27_valid_sink_size;
  reg [32-1:0] __reduce_max_27_valid_sink_stride;
  reg [32-1:0] __reduce_max_27_valid_sink_offset_buf;
  reg [33-1:0] __reduce_max_27_valid_sink_size_buf;
  reg [32-1:0] __reduce_max_27_valid_sink_stride_buf;
  reg [8-1:0] __reduce_max_27_valid_sink_sel;
  reg [32-1:0] __reduce_max_27_valid_sink_waddr;
  reg __reduce_max_27_valid_sink_wenable;
  reg [1-1:0] __reduce_max_27_valid_sink_wdata;
  reg __reduce_max_27_valid_sink_fifo_enq;
  reg [1-1:0] __reduce_max_27_valid_sink_fifo_wdata;
  reg [1-1:0] __reduce_max_27_valid_sink_immediate;
  reg _stream_conv2d_4_stream_ivalid;
  wire _stream_conv2d_4_stream_oready;
  wire _stream_conv2d_4_stream_internal_oready;
  assign _stream_conv2d_4_stream_oready = _stream_conv2d_4_stream_internal_oready;
  reg [32-1:0] _stream_conv2d_4_fsm;
  localparam _stream_conv2d_4_fsm_init = 0;
  wire _stream_conv2d_4_run_flag;
  reg _stream_conv2d_4_source_start;
  wire _stream_conv2d_4_source_stop;
  reg _stream_conv2d_4_source_busy;
  wire _stream_conv2d_4_sink_start;
  wire _stream_conv2d_4_sink_stop;
  wire _stream_conv2d_4_sink_busy;
  wire _stream_conv2d_4_busy;
  reg _stream_conv2d_4_busy_reg;
  wire _stream_conv2d_4_is_root;
  assign _stream_conv2d_4_is_root = 1;
  reg [1-1:0] _stream_conv2d_4_parameter_0_next_parameter_data;
  reg [2-1:0] _stream_conv2d_4_parameter_1_next_parameter_data;
  reg [2-1:0] _stream_conv2d_4_parameter_2_next_parameter_data;
  reg [9-1:0] _stream_conv2d_4_parameter_3_next_parameter_data;
  reg [1-1:0] _stream_conv2d_4_parameter_4_next_parameter_data;
  reg [1-1:0] _stream_conv2d_4_parameter_6_next_parameter_data;
  reg _stream_conv2d_4_source_7_idle;
  reg [33-1:0] _stream_conv2d_4_source_7_source_count;
  reg [5-1:0] _stream_conv2d_4_source_7_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_7_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_7_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_7_source_size;
  reg [32-1:0] _stream_conv2d_4_source_7_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_7_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_7_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_7_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_7_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_7_source_ram_raddr;
  reg _stream_conv2d_4_source_7_source_ram_renable;
  wire [16-1:0] _stream_conv2d_4_source_7_source_ram_rdata;
  reg _stream_conv2d_4_source_7_source_fifo_deq;
  wire [16-1:0] _stream_conv2d_4_source_7_source_fifo_rdata;
  reg [16-1:0] _stream_conv2d_4_source_7_source_empty_data;
  reg [1-1:0] _stream_conv2d_4_parameter_8_next_parameter_data;
  reg _stream_conv2d_4_source_9_idle;
  reg [33-1:0] _stream_conv2d_4_source_9_source_count;
  reg [5-1:0] _stream_conv2d_4_source_9_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_9_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_9_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_9_source_size;
  reg [32-1:0] _stream_conv2d_4_source_9_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_9_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_9_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_9_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_9_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_9_source_ram_raddr;
  reg _stream_conv2d_4_source_9_source_ram_renable;
  wire [16-1:0] _stream_conv2d_4_source_9_source_ram_rdata;
  reg _stream_conv2d_4_source_9_source_fifo_deq;
  wire [16-1:0] _stream_conv2d_4_source_9_source_fifo_rdata;
  reg [16-1:0] _stream_conv2d_4_source_9_source_empty_data;
  reg [1-1:0] _stream_conv2d_4_parameter_10_next_parameter_data;
  reg _stream_conv2d_4_source_11_idle;
  reg [33-1:0] _stream_conv2d_4_source_11_source_count;
  reg [5-1:0] _stream_conv2d_4_source_11_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_11_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_11_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_11_source_size;
  reg [32-1:0] _stream_conv2d_4_source_11_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_11_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_11_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_11_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_11_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_11_source_ram_raddr;
  reg _stream_conv2d_4_source_11_source_ram_renable;
  wire [16-1:0] _stream_conv2d_4_source_11_source_ram_rdata;
  reg _stream_conv2d_4_source_11_source_fifo_deq;
  wire [16-1:0] _stream_conv2d_4_source_11_source_fifo_rdata;
  reg [16-1:0] _stream_conv2d_4_source_11_source_empty_data;
  reg [1-1:0] _stream_conv2d_4_parameter_12_next_parameter_data;
  reg _stream_conv2d_4_source_13_idle;
  reg [33-1:0] _stream_conv2d_4_source_13_source_count;
  reg [5-1:0] _stream_conv2d_4_source_13_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_13_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_13_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_13_source_size;
  reg [32-1:0] _stream_conv2d_4_source_13_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_13_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_13_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_13_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_13_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_13_source_ram_raddr;
  reg _stream_conv2d_4_source_13_source_ram_renable;
  wire [16-1:0] _stream_conv2d_4_source_13_source_ram_rdata;
  reg _stream_conv2d_4_source_13_source_fifo_deq;
  wire [16-1:0] _stream_conv2d_4_source_13_source_fifo_rdata;
  reg [16-1:0] _stream_conv2d_4_source_13_source_empty_data;
  reg [1-1:0] _stream_conv2d_4_parameter_14_next_parameter_data;
  reg _stream_conv2d_4_source_15_idle;
  reg [33-1:0] _stream_conv2d_4_source_15_source_count;
  reg [5-1:0] _stream_conv2d_4_source_15_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_15_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_15_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_15_source_size;
  reg [32-1:0] _stream_conv2d_4_source_15_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_15_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_15_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_15_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_15_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_15_source_ram_raddr;
  reg _stream_conv2d_4_source_15_source_ram_renable;
  wire [16-1:0] _stream_conv2d_4_source_15_source_ram_rdata;
  reg _stream_conv2d_4_source_15_source_fifo_deq;
  wire [16-1:0] _stream_conv2d_4_source_15_source_fifo_rdata;
  reg [16-1:0] _stream_conv2d_4_source_15_source_empty_data;
  reg [1-1:0] _stream_conv2d_4_parameter_16_next_parameter_data;
  reg [1-1:0] _stream_conv2d_4_parameter_17_next_parameter_data;
  reg [5-1:0] _stream_conv2d_4_parameter_18_next_parameter_data;
  reg [1-1:0] _stream_conv2d_4_parameter_19_next_parameter_data;
  reg _stream_conv2d_4_source_20_idle;
  reg [33-1:0] _stream_conv2d_4_source_20_source_count;
  reg [5-1:0] _stream_conv2d_4_source_20_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_20_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_20_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_20_source_size;
  reg [32-1:0] _stream_conv2d_4_source_20_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_20_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_20_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_20_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_20_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_20_source_ram_raddr;
  reg _stream_conv2d_4_source_20_source_ram_renable;
  wire [16-1:0] _stream_conv2d_4_source_20_source_ram_rdata;
  reg _stream_conv2d_4_source_20_source_fifo_deq;
  wire [16-1:0] _stream_conv2d_4_source_20_source_fifo_rdata;
  reg [16-1:0] _stream_conv2d_4_source_20_source_empty_data;
  reg _stream_conv2d_4_source_21_idle;
  reg [33-1:0] _stream_conv2d_4_source_21_source_count;
  reg [5-1:0] _stream_conv2d_4_source_21_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_21_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_21_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_21_source_size;
  reg [32-1:0] _stream_conv2d_4_source_21_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_21_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_21_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_21_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_21_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_21_source_ram_raddr;
  reg _stream_conv2d_4_source_21_source_ram_renable;
  wire [16-1:0] _stream_conv2d_4_source_21_source_ram_rdata;
  reg _stream_conv2d_4_source_21_source_fifo_deq;
  wire [16-1:0] _stream_conv2d_4_source_21_source_fifo_rdata;
  reg [16-1:0] _stream_conv2d_4_source_21_source_empty_data;
  reg _stream_conv2d_4_source_22_idle;
  reg [33-1:0] _stream_conv2d_4_source_22_source_count;
  reg [5-1:0] _stream_conv2d_4_source_22_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_22_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_22_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_22_source_size;
  reg [32-1:0] _stream_conv2d_4_source_22_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_22_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_22_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_22_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_22_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_22_source_ram_raddr;
  reg _stream_conv2d_4_source_22_source_ram_renable;
  wire [16-1:0] _stream_conv2d_4_source_22_source_ram_rdata;
  reg _stream_conv2d_4_source_22_source_fifo_deq;
  wire [16-1:0] _stream_conv2d_4_source_22_source_fifo_rdata;
  reg [16-1:0] _stream_conv2d_4_source_22_source_empty_data;
  reg _stream_conv2d_4_source_23_idle;
  reg [33-1:0] _stream_conv2d_4_source_23_source_count;
  reg [5-1:0] _stream_conv2d_4_source_23_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_23_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_23_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_23_source_size;
  reg [32-1:0] _stream_conv2d_4_source_23_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_23_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_23_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_23_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_23_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_23_source_ram_raddr;
  reg _stream_conv2d_4_source_23_source_ram_renable;
  wire [16-1:0] _stream_conv2d_4_source_23_source_ram_rdata;
  reg _stream_conv2d_4_source_23_source_fifo_deq;
  wire [16-1:0] _stream_conv2d_4_source_23_source_fifo_rdata;
  reg [16-1:0] _stream_conv2d_4_source_23_source_empty_data;
  reg _stream_conv2d_4_source_24_idle;
  reg [33-1:0] _stream_conv2d_4_source_24_source_count;
  reg [5-1:0] _stream_conv2d_4_source_24_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_24_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_24_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_24_source_size;
  reg [32-1:0] _stream_conv2d_4_source_24_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_24_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_24_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_24_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_24_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_24_source_ram_raddr;
  reg _stream_conv2d_4_source_24_source_ram_renable;
  wire [16-1:0] _stream_conv2d_4_source_24_source_ram_rdata;
  reg _stream_conv2d_4_source_24_source_fifo_deq;
  wire [16-1:0] _stream_conv2d_4_source_24_source_fifo_rdata;
  reg [16-1:0] _stream_conv2d_4_source_24_source_empty_data;
  reg _stream_conv2d_4_source_25_idle;
  reg [33-1:0] _stream_conv2d_4_source_25_source_count;
  reg [5-1:0] _stream_conv2d_4_source_25_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_25_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_25_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_25_source_size;
  reg [32-1:0] _stream_conv2d_4_source_25_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_25_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_25_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_25_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_25_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_25_source_ram_raddr;
  reg _stream_conv2d_4_source_25_source_ram_renable;
  wire [16-1:0] _stream_conv2d_4_source_25_source_ram_rdata;
  reg _stream_conv2d_4_source_25_source_fifo_deq;
  wire [16-1:0] _stream_conv2d_4_source_25_source_fifo_rdata;
  reg [16-1:0] _stream_conv2d_4_source_25_source_empty_data;
  reg _stream_conv2d_4_source_26_idle;
  reg [33-1:0] _stream_conv2d_4_source_26_source_count;
  reg [5-1:0] _stream_conv2d_4_source_26_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_26_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_26_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_26_source_size;
  reg [32-1:0] _stream_conv2d_4_source_26_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_26_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_26_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_26_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_26_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_26_source_ram_raddr;
  reg _stream_conv2d_4_source_26_source_ram_renable;
  wire [16-1:0] _stream_conv2d_4_source_26_source_ram_rdata;
  reg _stream_conv2d_4_source_26_source_fifo_deq;
  wire [16-1:0] _stream_conv2d_4_source_26_source_fifo_rdata;
  reg [16-1:0] _stream_conv2d_4_source_26_source_empty_data;
  reg _stream_conv2d_4_source_27_idle;
  reg [33-1:0] _stream_conv2d_4_source_27_source_count;
  reg [5-1:0] _stream_conv2d_4_source_27_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_27_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_27_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_27_source_size;
  reg [32-1:0] _stream_conv2d_4_source_27_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_27_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_27_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_27_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_27_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_27_source_ram_raddr;
  reg _stream_conv2d_4_source_27_source_ram_renable;
  wire [16-1:0] _stream_conv2d_4_source_27_source_ram_rdata;
  reg _stream_conv2d_4_source_27_source_fifo_deq;
  wire [16-1:0] _stream_conv2d_4_source_27_source_fifo_rdata;
  reg [16-1:0] _stream_conv2d_4_source_27_source_empty_data;
  reg _stream_conv2d_4_source_28_idle;
  reg [33-1:0] _stream_conv2d_4_source_28_source_count;
  reg [5-1:0] _stream_conv2d_4_source_28_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_28_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_28_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_28_source_size;
  reg [32-1:0] _stream_conv2d_4_source_28_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_28_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_28_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_28_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_28_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_28_source_ram_raddr;
  reg _stream_conv2d_4_source_28_source_ram_renable;
  wire [16-1:0] _stream_conv2d_4_source_28_source_ram_rdata;
  reg _stream_conv2d_4_source_28_source_fifo_deq;
  wire [16-1:0] _stream_conv2d_4_source_28_source_fifo_rdata;
  reg [16-1:0] _stream_conv2d_4_source_28_source_empty_data;
  reg _stream_conv2d_4_source_29_idle;
  reg [33-1:0] _stream_conv2d_4_source_29_source_count;
  reg [5-1:0] _stream_conv2d_4_source_29_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_29_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_29_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_29_source_size;
  reg [32-1:0] _stream_conv2d_4_source_29_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_29_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_29_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_29_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_29_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_29_source_ram_raddr;
  reg _stream_conv2d_4_source_29_source_ram_renable;
  wire [16-1:0] _stream_conv2d_4_source_29_source_ram_rdata;
  reg _stream_conv2d_4_source_29_source_fifo_deq;
  wire [16-1:0] _stream_conv2d_4_source_29_source_fifo_rdata;
  reg [16-1:0] _stream_conv2d_4_source_29_source_empty_data;
  reg _stream_conv2d_4_source_30_idle;
  reg [33-1:0] _stream_conv2d_4_source_30_source_count;
  reg [5-1:0] _stream_conv2d_4_source_30_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_30_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_30_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_30_source_size;
  reg [32-1:0] _stream_conv2d_4_source_30_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_30_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_30_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_30_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_30_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_30_source_ram_raddr;
  reg _stream_conv2d_4_source_30_source_ram_renable;
  wire [16-1:0] _stream_conv2d_4_source_30_source_ram_rdata;
  reg _stream_conv2d_4_source_30_source_fifo_deq;
  wire [16-1:0] _stream_conv2d_4_source_30_source_fifo_rdata;
  reg [16-1:0] _stream_conv2d_4_source_30_source_empty_data;
  reg _stream_conv2d_4_source_31_idle;
  reg [33-1:0] _stream_conv2d_4_source_31_source_count;
  reg [5-1:0] _stream_conv2d_4_source_31_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_31_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_31_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_31_source_size;
  reg [32-1:0] _stream_conv2d_4_source_31_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_31_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_31_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_31_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_31_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_31_source_ram_raddr;
  reg _stream_conv2d_4_source_31_source_ram_renable;
  wire [16-1:0] _stream_conv2d_4_source_31_source_ram_rdata;
  reg _stream_conv2d_4_source_31_source_fifo_deq;
  wire [16-1:0] _stream_conv2d_4_source_31_source_fifo_rdata;
  reg [16-1:0] _stream_conv2d_4_source_31_source_empty_data;
  reg _stream_conv2d_4_source_32_idle;
  reg [33-1:0] _stream_conv2d_4_source_32_source_count;
  reg [5-1:0] _stream_conv2d_4_source_32_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_32_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_32_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_32_source_size;
  reg [32-1:0] _stream_conv2d_4_source_32_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_32_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_32_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_32_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_32_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_32_source_ram_raddr;
  reg _stream_conv2d_4_source_32_source_ram_renable;
  wire [16-1:0] _stream_conv2d_4_source_32_source_ram_rdata;
  reg _stream_conv2d_4_source_32_source_fifo_deq;
  wire [16-1:0] _stream_conv2d_4_source_32_source_fifo_rdata;
  reg [16-1:0] _stream_conv2d_4_source_32_source_empty_data;
  reg _stream_conv2d_4_source_33_idle;
  reg [33-1:0] _stream_conv2d_4_source_33_source_count;
  reg [5-1:0] _stream_conv2d_4_source_33_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_33_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_33_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_33_source_size;
  reg [32-1:0] _stream_conv2d_4_source_33_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_33_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_33_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_33_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_33_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_33_source_ram_raddr;
  reg _stream_conv2d_4_source_33_source_ram_renable;
  wire [16-1:0] _stream_conv2d_4_source_33_source_ram_rdata;
  reg _stream_conv2d_4_source_33_source_fifo_deq;
  wire [16-1:0] _stream_conv2d_4_source_33_source_fifo_rdata;
  reg [16-1:0] _stream_conv2d_4_source_33_source_empty_data;
  reg _stream_conv2d_4_source_34_idle;
  reg [33-1:0] _stream_conv2d_4_source_34_source_count;
  reg [5-1:0] _stream_conv2d_4_source_34_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_34_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_34_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_34_source_size;
  reg [32-1:0] _stream_conv2d_4_source_34_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_34_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_34_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_34_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_34_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_34_source_ram_raddr;
  reg _stream_conv2d_4_source_34_source_ram_renable;
  wire [16-1:0] _stream_conv2d_4_source_34_source_ram_rdata;
  reg _stream_conv2d_4_source_34_source_fifo_deq;
  wire [16-1:0] _stream_conv2d_4_source_34_source_fifo_rdata;
  reg [16-1:0] _stream_conv2d_4_source_34_source_empty_data;
  reg _stream_conv2d_4_source_35_idle;
  reg [33-1:0] _stream_conv2d_4_source_35_source_count;
  reg [5-1:0] _stream_conv2d_4_source_35_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_35_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_35_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_35_source_size;
  reg [32-1:0] _stream_conv2d_4_source_35_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_35_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_35_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_35_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_35_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_35_source_ram_raddr;
  reg _stream_conv2d_4_source_35_source_ram_renable;
  wire [16-1:0] _stream_conv2d_4_source_35_source_ram_rdata;
  reg _stream_conv2d_4_source_35_source_fifo_deq;
  wire [16-1:0] _stream_conv2d_4_source_35_source_fifo_rdata;
  reg [16-1:0] _stream_conv2d_4_source_35_source_empty_data;
  reg _stream_conv2d_4_source_36_idle;
  reg [33-1:0] _stream_conv2d_4_source_36_source_count;
  reg [5-1:0] _stream_conv2d_4_source_36_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_36_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_36_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_36_source_size;
  reg [32-1:0] _stream_conv2d_4_source_36_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_36_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_36_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_36_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_36_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_36_source_ram_raddr;
  reg _stream_conv2d_4_source_36_source_ram_renable;
  wire [16-1:0] _stream_conv2d_4_source_36_source_ram_rdata;
  reg _stream_conv2d_4_source_36_source_fifo_deq;
  wire [16-1:0] _stream_conv2d_4_source_36_source_fifo_rdata;
  reg [16-1:0] _stream_conv2d_4_source_36_source_empty_data;
  reg _stream_conv2d_4_source_37_idle;
  reg [33-1:0] _stream_conv2d_4_source_37_source_count;
  reg [5-1:0] _stream_conv2d_4_source_37_source_mode;
  reg [16-1:0] _stream_conv2d_4_source_37_source_generator_id;
  reg [32-1:0] _stream_conv2d_4_source_37_source_offset;
  reg [33-1:0] _stream_conv2d_4_source_37_source_size;
  reg [32-1:0] _stream_conv2d_4_source_37_source_stride;
  reg [32-1:0] _stream_conv2d_4_source_37_source_offset_buf;
  reg [33-1:0] _stream_conv2d_4_source_37_source_size_buf;
  reg [32-1:0] _stream_conv2d_4_source_37_source_stride_buf;
  reg [8-1:0] _stream_conv2d_4_source_37_source_sel;
  reg [32-1:0] _stream_conv2d_4_source_37_source_ram_raddr;
  reg _stream_conv2d_4_source_37_source_ram_renable;
  wire [16-1:0] _stream_conv2d_4_source_37_source_ram_rdata;
  reg _stream_conv2d_4_source_37_source_fifo_deq;
  wire [16-1:0] _stream_conv2d_4_source_37_source_fifo_rdata;
  reg [16-1:0] _stream_conv2d_4_source_37_source_empty_data;
  wire signed [16-1:0] mul_18_x_data;
  wire signed [16-1:0] mul_18_y_data;
  wire [5-1:0] mul_18_rshift_data;
  reg __mul_18_stream_ivalid_1;
  reg __mul_18_stream_ivalid_2;
  reg __mul_18_stream_ivalid_3;
  reg __mul_18_stream_ivalid_4;
  reg __mul_18_stream_ivalid_5;
  reg __mul_18_stream_ivalid_6;
  reg __mul_18_stream_ivalid_7;
  reg __mul_18_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_1355;
  reg [5-1:0] _minus_data_1357;
  reg [1-1:0] _greatereq_data_1368;
  reg signed [16-1:0] __delay_data_1930__variable_1352;
  reg signed [16-1:0] __delay_data_1933__variable_1353;
  reg [5-1:0] __delay_data_1936__variable_1354;
  reg signed [34-1:0] _sll_data_1359;
  reg [1-1:0] __delay_data_1927_greaterthan_1355;
  reg [1-1:0] __delay_data_1928_greatereq_1368;
  reg signed [16-1:0] __delay_data_1931__delay_1930__variable_1352;
  reg signed [16-1:0] __delay_data_1934__delay_1933__variable_1353;
  reg [5-1:0] __delay_data_1937__delay_1936__variable_1354;
  reg signed [32-1:0] _cond_data_1365;
  reg [1-1:0] __delay_data_1929__delay_1928_greatereq_1368;
  reg signed [16-1:0] __delay_data_1932__delay_1931__delay_1930__variable_1352;
  reg signed [16-1:0] __delay_data_1935__delay_1934__delay_1933__variable_1353;
  reg [5-1:0] __delay_data_1938__delay_1937__delay_1936__variable_1354;
  wire signed [16-1:0] _uminus_data_1367;
  assign _uminus_data_1367 = -_cond_data_1365;
  wire signed [16-1:0] _cond_data_1370;
  assign _cond_data_1370 = (__delay_data_1929__delay_1928_greatereq_1368)? _cond_data_1365 : _uminus_data_1367;
  wire signed [32-1:0] __muladd_madd_odata_1371;
  reg signed [32-1:0] __muladd_madd_odata_reg_1371;
  wire signed [32-1:0] __muladd_data_1371;
  assign __muladd_data_1371 = __muladd_madd_odata_reg_1371;
  wire __muladd_madd_update_1371;
  assign __muladd_madd_update_1371 = _mul_18_stream_oready;

  madd_9
  __muladd_madd_1371
  (
    .CLK(CLK),
    .update(__muladd_madd_update_1371),
    .a(__delay_data_1932__delay_1931__delay_1930__variable_1352),
    .b(__delay_data_1935__delay_1934__delay_1933__variable_1353),
    .c(_cond_data_1370),
    .d(__muladd_madd_odata_1371)
  );

  reg [5-1:0] __delay_data_1939__delay_1938__delay_1937____variable_1354;
  reg [5-1:0] __delay_data_1940__delay_1939__delay_1938____variable_1354;
  reg [5-1:0] __delay_data_1941__delay_1940__delay_1939____variable_1354;
  reg [5-1:0] __delay_data_1942__delay_1941__delay_1940____variable_1354;
  reg signed [32-1:0] _sra_data_1372;
  wire signed [32-1:0] mul_18_z_data;
  assign mul_18_z_data = _sra_data_1372;
  wire signed [16-1:0] mul_19_x_data;
  wire signed [16-1:0] mul_19_y_data;
  wire [5-1:0] mul_19_rshift_data;
  reg __mul_19_stream_ivalid_1;
  reg __mul_19_stream_ivalid_2;
  reg __mul_19_stream_ivalid_3;
  reg __mul_19_stream_ivalid_4;
  reg __mul_19_stream_ivalid_5;
  reg __mul_19_stream_ivalid_6;
  reg __mul_19_stream_ivalid_7;
  reg __mul_19_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_1376;
  reg [5-1:0] _minus_data_1378;
  reg [1-1:0] _greatereq_data_1389;
  reg signed [16-1:0] __delay_data_1949__variable_1373;
  reg signed [16-1:0] __delay_data_1952__variable_1374;
  reg [5-1:0] __delay_data_1955__variable_1375;
  reg signed [34-1:0] _sll_data_1380;
  reg [1-1:0] __delay_data_1946_greaterthan_1376;
  reg [1-1:0] __delay_data_1947_greatereq_1389;
  reg signed [16-1:0] __delay_data_1950__delay_1949__variable_1373;
  reg signed [16-1:0] __delay_data_1953__delay_1952__variable_1374;
  reg [5-1:0] __delay_data_1956__delay_1955__variable_1375;
  reg signed [32-1:0] _cond_data_1386;
  reg [1-1:0] __delay_data_1948__delay_1947_greatereq_1389;
  reg signed [16-1:0] __delay_data_1951__delay_1950__delay_1949__variable_1373;
  reg signed [16-1:0] __delay_data_1954__delay_1953__delay_1952__variable_1374;
  reg [5-1:0] __delay_data_1957__delay_1956__delay_1955__variable_1375;
  wire signed [16-1:0] _uminus_data_1388;
  assign _uminus_data_1388 = -_cond_data_1386;
  wire signed [16-1:0] _cond_data_1391;
  assign _cond_data_1391 = (__delay_data_1948__delay_1947_greatereq_1389)? _cond_data_1386 : _uminus_data_1388;
  wire signed [32-1:0] __muladd_madd_odata_1392;
  reg signed [32-1:0] __muladd_madd_odata_reg_1392;
  wire signed [32-1:0] __muladd_data_1392;
  assign __muladd_data_1392 = __muladd_madd_odata_reg_1392;
  wire __muladd_madd_update_1392;
  assign __muladd_madd_update_1392 = _mul_19_stream_oready;

  madd_10
  __muladd_madd_1392
  (
    .CLK(CLK),
    .update(__muladd_madd_update_1392),
    .a(__delay_data_1951__delay_1950__delay_1949__variable_1373),
    .b(__delay_data_1954__delay_1953__delay_1952__variable_1374),
    .c(_cond_data_1391),
    .d(__muladd_madd_odata_1392)
  );

  reg [5-1:0] __delay_data_1958__delay_1957__delay_1956____variable_1375;
  reg [5-1:0] __delay_data_1959__delay_1958__delay_1957____variable_1375;
  reg [5-1:0] __delay_data_1960__delay_1959__delay_1958____variable_1375;
  reg [5-1:0] __delay_data_1961__delay_1960__delay_1959____variable_1375;
  reg signed [32-1:0] _sra_data_1393;
  wire signed [32-1:0] mul_19_z_data;
  assign mul_19_z_data = _sra_data_1393;
  wire signed [16-1:0] mul_20_x_data;
  wire signed [16-1:0] mul_20_y_data;
  wire [5-1:0] mul_20_rshift_data;
  reg __mul_20_stream_ivalid_1;
  reg __mul_20_stream_ivalid_2;
  reg __mul_20_stream_ivalid_3;
  reg __mul_20_stream_ivalid_4;
  reg __mul_20_stream_ivalid_5;
  reg __mul_20_stream_ivalid_6;
  reg __mul_20_stream_ivalid_7;
  reg __mul_20_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_1397;
  reg [5-1:0] _minus_data_1399;
  reg [1-1:0] _greatereq_data_1410;
  reg signed [16-1:0] __delay_data_1968__variable_1394;
  reg signed [16-1:0] __delay_data_1971__variable_1395;
  reg [5-1:0] __delay_data_1974__variable_1396;
  reg signed [34-1:0] _sll_data_1401;
  reg [1-1:0] __delay_data_1965_greaterthan_1397;
  reg [1-1:0] __delay_data_1966_greatereq_1410;
  reg signed [16-1:0] __delay_data_1969__delay_1968__variable_1394;
  reg signed [16-1:0] __delay_data_1972__delay_1971__variable_1395;
  reg [5-1:0] __delay_data_1975__delay_1974__variable_1396;
  reg signed [32-1:0] _cond_data_1407;
  reg [1-1:0] __delay_data_1967__delay_1966_greatereq_1410;
  reg signed [16-1:0] __delay_data_1970__delay_1969__delay_1968__variable_1394;
  reg signed [16-1:0] __delay_data_1973__delay_1972__delay_1971__variable_1395;
  reg [5-1:0] __delay_data_1976__delay_1975__delay_1974__variable_1396;
  wire signed [16-1:0] _uminus_data_1409;
  assign _uminus_data_1409 = -_cond_data_1407;
  wire signed [16-1:0] _cond_data_1412;
  assign _cond_data_1412 = (__delay_data_1967__delay_1966_greatereq_1410)? _cond_data_1407 : _uminus_data_1409;
  wire signed [32-1:0] __muladd_madd_odata_1413;
  reg signed [32-1:0] __muladd_madd_odata_reg_1413;
  wire signed [32-1:0] __muladd_data_1413;
  assign __muladd_data_1413 = __muladd_madd_odata_reg_1413;
  wire __muladd_madd_update_1413;
  assign __muladd_madd_update_1413 = _mul_20_stream_oready;

  madd_11
  __muladd_madd_1413
  (
    .CLK(CLK),
    .update(__muladd_madd_update_1413),
    .a(__delay_data_1970__delay_1969__delay_1968__variable_1394),
    .b(__delay_data_1973__delay_1972__delay_1971__variable_1395),
    .c(_cond_data_1412),
    .d(__muladd_madd_odata_1413)
  );

  reg [5-1:0] __delay_data_1977__delay_1976__delay_1975____variable_1396;
  reg [5-1:0] __delay_data_1978__delay_1977__delay_1976____variable_1396;
  reg [5-1:0] __delay_data_1979__delay_1978__delay_1977____variable_1396;
  reg [5-1:0] __delay_data_1980__delay_1979__delay_1978____variable_1396;
  reg signed [32-1:0] _sra_data_1414;
  wire signed [32-1:0] mul_20_z_data;
  assign mul_20_z_data = _sra_data_1414;
  wire signed [16-1:0] mul_21_x_data;
  wire signed [16-1:0] mul_21_y_data;
  wire [5-1:0] mul_21_rshift_data;
  reg __mul_21_stream_ivalid_1;
  reg __mul_21_stream_ivalid_2;
  reg __mul_21_stream_ivalid_3;
  reg __mul_21_stream_ivalid_4;
  reg __mul_21_stream_ivalid_5;
  reg __mul_21_stream_ivalid_6;
  reg __mul_21_stream_ivalid_7;
  reg __mul_21_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_1418;
  reg [5-1:0] _minus_data_1420;
  reg [1-1:0] _greatereq_data_1431;
  reg signed [16-1:0] __delay_data_1987__variable_1415;
  reg signed [16-1:0] __delay_data_1990__variable_1416;
  reg [5-1:0] __delay_data_1993__variable_1417;
  reg signed [34-1:0] _sll_data_1422;
  reg [1-1:0] __delay_data_1984_greaterthan_1418;
  reg [1-1:0] __delay_data_1985_greatereq_1431;
  reg signed [16-1:0] __delay_data_1988__delay_1987__variable_1415;
  reg signed [16-1:0] __delay_data_1991__delay_1990__variable_1416;
  reg [5-1:0] __delay_data_1994__delay_1993__variable_1417;
  reg signed [32-1:0] _cond_data_1428;
  reg [1-1:0] __delay_data_1986__delay_1985_greatereq_1431;
  reg signed [16-1:0] __delay_data_1989__delay_1988__delay_1987__variable_1415;
  reg signed [16-1:0] __delay_data_1992__delay_1991__delay_1990__variable_1416;
  reg [5-1:0] __delay_data_1995__delay_1994__delay_1993__variable_1417;
  wire signed [16-1:0] _uminus_data_1430;
  assign _uminus_data_1430 = -_cond_data_1428;
  wire signed [16-1:0] _cond_data_1433;
  assign _cond_data_1433 = (__delay_data_1986__delay_1985_greatereq_1431)? _cond_data_1428 : _uminus_data_1430;
  wire signed [32-1:0] __muladd_madd_odata_1434;
  reg signed [32-1:0] __muladd_madd_odata_reg_1434;
  wire signed [32-1:0] __muladd_data_1434;
  assign __muladd_data_1434 = __muladd_madd_odata_reg_1434;
  wire __muladd_madd_update_1434;
  assign __muladd_madd_update_1434 = _mul_21_stream_oready;

  madd_12
  __muladd_madd_1434
  (
    .CLK(CLK),
    .update(__muladd_madd_update_1434),
    .a(__delay_data_1989__delay_1988__delay_1987__variable_1415),
    .b(__delay_data_1992__delay_1991__delay_1990__variable_1416),
    .c(_cond_data_1433),
    .d(__muladd_madd_odata_1434)
  );

  reg [5-1:0] __delay_data_1996__delay_1995__delay_1994____variable_1417;
  reg [5-1:0] __delay_data_1997__delay_1996__delay_1995____variable_1417;
  reg [5-1:0] __delay_data_1998__delay_1997__delay_1996____variable_1417;
  reg [5-1:0] __delay_data_1999__delay_1998__delay_1997____variable_1417;
  reg signed [32-1:0] _sra_data_1435;
  wire signed [32-1:0] mul_21_z_data;
  assign mul_21_z_data = _sra_data_1435;
  wire signed [16-1:0] mul_22_x_data;
  wire signed [16-1:0] mul_22_y_data;
  wire [5-1:0] mul_22_rshift_data;
  reg __mul_22_stream_ivalid_1;
  reg __mul_22_stream_ivalid_2;
  reg __mul_22_stream_ivalid_3;
  reg __mul_22_stream_ivalid_4;
  reg __mul_22_stream_ivalid_5;
  reg __mul_22_stream_ivalid_6;
  reg __mul_22_stream_ivalid_7;
  reg __mul_22_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_1439;
  reg [5-1:0] _minus_data_1441;
  reg [1-1:0] _greatereq_data_1452;
  reg signed [16-1:0] __delay_data_2006__variable_1436;
  reg signed [16-1:0] __delay_data_2009__variable_1437;
  reg [5-1:0] __delay_data_2012__variable_1438;
  reg signed [34-1:0] _sll_data_1443;
  reg [1-1:0] __delay_data_2003_greaterthan_1439;
  reg [1-1:0] __delay_data_2004_greatereq_1452;
  reg signed [16-1:0] __delay_data_2007__delay_2006__variable_1436;
  reg signed [16-1:0] __delay_data_2010__delay_2009__variable_1437;
  reg [5-1:0] __delay_data_2013__delay_2012__variable_1438;
  reg signed [32-1:0] _cond_data_1449;
  reg [1-1:0] __delay_data_2005__delay_2004_greatereq_1452;
  reg signed [16-1:0] __delay_data_2008__delay_2007__delay_2006__variable_1436;
  reg signed [16-1:0] __delay_data_2011__delay_2010__delay_2009__variable_1437;
  reg [5-1:0] __delay_data_2014__delay_2013__delay_2012__variable_1438;
  wire signed [16-1:0] _uminus_data_1451;
  assign _uminus_data_1451 = -_cond_data_1449;
  wire signed [16-1:0] _cond_data_1454;
  assign _cond_data_1454 = (__delay_data_2005__delay_2004_greatereq_1452)? _cond_data_1449 : _uminus_data_1451;
  wire signed [32-1:0] __muladd_madd_odata_1455;
  reg signed [32-1:0] __muladd_madd_odata_reg_1455;
  wire signed [32-1:0] __muladd_data_1455;
  assign __muladd_data_1455 = __muladd_madd_odata_reg_1455;
  wire __muladd_madd_update_1455;
  assign __muladd_madd_update_1455 = _mul_22_stream_oready;

  madd_13
  __muladd_madd_1455
  (
    .CLK(CLK),
    .update(__muladd_madd_update_1455),
    .a(__delay_data_2008__delay_2007__delay_2006__variable_1436),
    .b(__delay_data_2011__delay_2010__delay_2009__variable_1437),
    .c(_cond_data_1454),
    .d(__muladd_madd_odata_1455)
  );

  reg [5-1:0] __delay_data_2015__delay_2014__delay_2013____variable_1438;
  reg [5-1:0] __delay_data_2016__delay_2015__delay_2014____variable_1438;
  reg [5-1:0] __delay_data_2017__delay_2016__delay_2015____variable_1438;
  reg [5-1:0] __delay_data_2018__delay_2017__delay_2016____variable_1438;
  reg signed [32-1:0] _sra_data_1456;
  wire signed [32-1:0] mul_22_z_data;
  assign mul_22_z_data = _sra_data_1456;
  wire signed [16-1:0] mul_23_x_data;
  wire signed [16-1:0] mul_23_y_data;
  wire [5-1:0] mul_23_rshift_data;
  reg __mul_23_stream_ivalid_1;
  reg __mul_23_stream_ivalid_2;
  reg __mul_23_stream_ivalid_3;
  reg __mul_23_stream_ivalid_4;
  reg __mul_23_stream_ivalid_5;
  reg __mul_23_stream_ivalid_6;
  reg __mul_23_stream_ivalid_7;
  reg __mul_23_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_1460;
  reg [5-1:0] _minus_data_1462;
  reg [1-1:0] _greatereq_data_1473;
  reg signed [16-1:0] __delay_data_2025__variable_1457;
  reg signed [16-1:0] __delay_data_2028__variable_1458;
  reg [5-1:0] __delay_data_2031__variable_1459;
  reg signed [34-1:0] _sll_data_1464;
  reg [1-1:0] __delay_data_2022_greaterthan_1460;
  reg [1-1:0] __delay_data_2023_greatereq_1473;
  reg signed [16-1:0] __delay_data_2026__delay_2025__variable_1457;
  reg signed [16-1:0] __delay_data_2029__delay_2028__variable_1458;
  reg [5-1:0] __delay_data_2032__delay_2031__variable_1459;
  reg signed [32-1:0] _cond_data_1470;
  reg [1-1:0] __delay_data_2024__delay_2023_greatereq_1473;
  reg signed [16-1:0] __delay_data_2027__delay_2026__delay_2025__variable_1457;
  reg signed [16-1:0] __delay_data_2030__delay_2029__delay_2028__variable_1458;
  reg [5-1:0] __delay_data_2033__delay_2032__delay_2031__variable_1459;
  wire signed [16-1:0] _uminus_data_1472;
  assign _uminus_data_1472 = -_cond_data_1470;
  wire signed [16-1:0] _cond_data_1475;
  assign _cond_data_1475 = (__delay_data_2024__delay_2023_greatereq_1473)? _cond_data_1470 : _uminus_data_1472;
  wire signed [32-1:0] __muladd_madd_odata_1476;
  reg signed [32-1:0] __muladd_madd_odata_reg_1476;
  wire signed [32-1:0] __muladd_data_1476;
  assign __muladd_data_1476 = __muladd_madd_odata_reg_1476;
  wire __muladd_madd_update_1476;
  assign __muladd_madd_update_1476 = _mul_23_stream_oready;

  madd_14
  __muladd_madd_1476
  (
    .CLK(CLK),
    .update(__muladd_madd_update_1476),
    .a(__delay_data_2027__delay_2026__delay_2025__variable_1457),
    .b(__delay_data_2030__delay_2029__delay_2028__variable_1458),
    .c(_cond_data_1475),
    .d(__muladd_madd_odata_1476)
  );

  reg [5-1:0] __delay_data_2034__delay_2033__delay_2032____variable_1459;
  reg [5-1:0] __delay_data_2035__delay_2034__delay_2033____variable_1459;
  reg [5-1:0] __delay_data_2036__delay_2035__delay_2034____variable_1459;
  reg [5-1:0] __delay_data_2037__delay_2036__delay_2035____variable_1459;
  reg signed [32-1:0] _sra_data_1477;
  wire signed [32-1:0] mul_23_z_data;
  assign mul_23_z_data = _sra_data_1477;
  wire signed [16-1:0] mul_24_x_data;
  wire signed [16-1:0] mul_24_y_data;
  wire [5-1:0] mul_24_rshift_data;
  reg __mul_24_stream_ivalid_1;
  reg __mul_24_stream_ivalid_2;
  reg __mul_24_stream_ivalid_3;
  reg __mul_24_stream_ivalid_4;
  reg __mul_24_stream_ivalid_5;
  reg __mul_24_stream_ivalid_6;
  reg __mul_24_stream_ivalid_7;
  reg __mul_24_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_1481;
  reg [5-1:0] _minus_data_1483;
  reg [1-1:0] _greatereq_data_1494;
  reg signed [16-1:0] __delay_data_2044__variable_1478;
  reg signed [16-1:0] __delay_data_2047__variable_1479;
  reg [5-1:0] __delay_data_2050__variable_1480;
  reg signed [34-1:0] _sll_data_1485;
  reg [1-1:0] __delay_data_2041_greaterthan_1481;
  reg [1-1:0] __delay_data_2042_greatereq_1494;
  reg signed [16-1:0] __delay_data_2045__delay_2044__variable_1478;
  reg signed [16-1:0] __delay_data_2048__delay_2047__variable_1479;
  reg [5-1:0] __delay_data_2051__delay_2050__variable_1480;
  reg signed [32-1:0] _cond_data_1491;
  reg [1-1:0] __delay_data_2043__delay_2042_greatereq_1494;
  reg signed [16-1:0] __delay_data_2046__delay_2045__delay_2044__variable_1478;
  reg signed [16-1:0] __delay_data_2049__delay_2048__delay_2047__variable_1479;
  reg [5-1:0] __delay_data_2052__delay_2051__delay_2050__variable_1480;
  wire signed [16-1:0] _uminus_data_1493;
  assign _uminus_data_1493 = -_cond_data_1491;
  wire signed [16-1:0] _cond_data_1496;
  assign _cond_data_1496 = (__delay_data_2043__delay_2042_greatereq_1494)? _cond_data_1491 : _uminus_data_1493;
  wire signed [32-1:0] __muladd_madd_odata_1497;
  reg signed [32-1:0] __muladd_madd_odata_reg_1497;
  wire signed [32-1:0] __muladd_data_1497;
  assign __muladd_data_1497 = __muladd_madd_odata_reg_1497;
  wire __muladd_madd_update_1497;
  assign __muladd_madd_update_1497 = _mul_24_stream_oready;

  madd_15
  __muladd_madd_1497
  (
    .CLK(CLK),
    .update(__muladd_madd_update_1497),
    .a(__delay_data_2046__delay_2045__delay_2044__variable_1478),
    .b(__delay_data_2049__delay_2048__delay_2047__variable_1479),
    .c(_cond_data_1496),
    .d(__muladd_madd_odata_1497)
  );

  reg [5-1:0] __delay_data_2053__delay_2052__delay_2051____variable_1480;
  reg [5-1:0] __delay_data_2054__delay_2053__delay_2052____variable_1480;
  reg [5-1:0] __delay_data_2055__delay_2054__delay_2053____variable_1480;
  reg [5-1:0] __delay_data_2056__delay_2055__delay_2054____variable_1480;
  reg signed [32-1:0] _sra_data_1498;
  wire signed [32-1:0] mul_24_z_data;
  assign mul_24_z_data = _sra_data_1498;
  wire signed [16-1:0] mul_25_x_data;
  wire signed [16-1:0] mul_25_y_data;
  wire [5-1:0] mul_25_rshift_data;
  reg __mul_25_stream_ivalid_1;
  reg __mul_25_stream_ivalid_2;
  reg __mul_25_stream_ivalid_3;
  reg __mul_25_stream_ivalid_4;
  reg __mul_25_stream_ivalid_5;
  reg __mul_25_stream_ivalid_6;
  reg __mul_25_stream_ivalid_7;
  reg __mul_25_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_1502;
  reg [5-1:0] _minus_data_1504;
  reg [1-1:0] _greatereq_data_1515;
  reg signed [16-1:0] __delay_data_2063__variable_1499;
  reg signed [16-1:0] __delay_data_2066__variable_1500;
  reg [5-1:0] __delay_data_2069__variable_1501;
  reg signed [34-1:0] _sll_data_1506;
  reg [1-1:0] __delay_data_2060_greaterthan_1502;
  reg [1-1:0] __delay_data_2061_greatereq_1515;
  reg signed [16-1:0] __delay_data_2064__delay_2063__variable_1499;
  reg signed [16-1:0] __delay_data_2067__delay_2066__variable_1500;
  reg [5-1:0] __delay_data_2070__delay_2069__variable_1501;
  reg signed [32-1:0] _cond_data_1512;
  reg [1-1:0] __delay_data_2062__delay_2061_greatereq_1515;
  reg signed [16-1:0] __delay_data_2065__delay_2064__delay_2063__variable_1499;
  reg signed [16-1:0] __delay_data_2068__delay_2067__delay_2066__variable_1500;
  reg [5-1:0] __delay_data_2071__delay_2070__delay_2069__variable_1501;
  wire signed [16-1:0] _uminus_data_1514;
  assign _uminus_data_1514 = -_cond_data_1512;
  wire signed [16-1:0] _cond_data_1517;
  assign _cond_data_1517 = (__delay_data_2062__delay_2061_greatereq_1515)? _cond_data_1512 : _uminus_data_1514;
  wire signed [32-1:0] __muladd_madd_odata_1518;
  reg signed [32-1:0] __muladd_madd_odata_reg_1518;
  wire signed [32-1:0] __muladd_data_1518;
  assign __muladd_data_1518 = __muladd_madd_odata_reg_1518;
  wire __muladd_madd_update_1518;
  assign __muladd_madd_update_1518 = _mul_25_stream_oready;

  madd_16
  __muladd_madd_1518
  (
    .CLK(CLK),
    .update(__muladd_madd_update_1518),
    .a(__delay_data_2065__delay_2064__delay_2063__variable_1499),
    .b(__delay_data_2068__delay_2067__delay_2066__variable_1500),
    .c(_cond_data_1517),
    .d(__muladd_madd_odata_1518)
  );

  reg [5-1:0] __delay_data_2072__delay_2071__delay_2070____variable_1501;
  reg [5-1:0] __delay_data_2073__delay_2072__delay_2071____variable_1501;
  reg [5-1:0] __delay_data_2074__delay_2073__delay_2072____variable_1501;
  reg [5-1:0] __delay_data_2075__delay_2074__delay_2073____variable_1501;
  reg signed [32-1:0] _sra_data_1519;
  wire signed [32-1:0] mul_25_z_data;
  assign mul_25_z_data = _sra_data_1519;
  wire signed [16-1:0] mul_26_x_data;
  wire signed [16-1:0] mul_26_y_data;
  wire [5-1:0] mul_26_rshift_data;
  reg __mul_26_stream_ivalid_1;
  reg __mul_26_stream_ivalid_2;
  reg __mul_26_stream_ivalid_3;
  reg __mul_26_stream_ivalid_4;
  reg __mul_26_stream_ivalid_5;
  reg __mul_26_stream_ivalid_6;
  reg __mul_26_stream_ivalid_7;
  reg __mul_26_stream_ivalid_8;
  reg [1-1:0] _greaterthan_data_1523;
  reg [5-1:0] _minus_data_1525;
  reg [1-1:0] _greatereq_data_1536;
  reg signed [16-1:0] __delay_data_2082__variable_1520;
  reg signed [16-1:0] __delay_data_2085__variable_1521;
  reg [5-1:0] __delay_data_2088__variable_1522;
  reg signed [34-1:0] _sll_data_1527;
  reg [1-1:0] __delay_data_2079_greaterthan_1523;
  reg [1-1:0] __delay_data_2080_greatereq_1536;
  reg signed [16-1:0] __delay_data_2083__delay_2082__variable_1520;
  reg signed [16-1:0] __delay_data_2086__delay_2085__variable_1521;
  reg [5-1:0] __delay_data_2089__delay_2088__variable_1522;
  reg signed [32-1:0] _cond_data_1533;
  reg [1-1:0] __delay_data_2081__delay_2080_greatereq_1536;
  reg signed [16-1:0] __delay_data_2084__delay_2083__delay_2082__variable_1520;
  reg signed [16-1:0] __delay_data_2087__delay_2086__delay_2085__variable_1521;
  reg [5-1:0] __delay_data_2090__delay_2089__delay_2088__variable_1522;
  wire signed [16-1:0] _uminus_data_1535;
  assign _uminus_data_1535 = -_cond_data_1533;
  wire signed [16-1:0] _cond_data_1538;
  assign _cond_data_1538 = (__delay_data_2081__delay_2080_greatereq_1536)? _cond_data_1533 : _uminus_data_1535;
  wire signed [32-1:0] __muladd_madd_odata_1539;
  reg signed [32-1:0] __muladd_madd_odata_reg_1539;
  wire signed [32-1:0] __muladd_data_1539;
  assign __muladd_data_1539 = __muladd_madd_odata_reg_1539;
  wire __muladd_madd_update_1539;
  assign __muladd_madd_update_1539 = _mul_26_stream_oready;

  madd_17
  __muladd_madd_1539
  (
    .CLK(CLK),
    .update(__muladd_madd_update_1539),
    .a(__delay_data_2084__delay_2083__delay_2082__variable_1520),
    .b(__delay_data_2087__delay_2086__delay_2085__variable_1521),
    .c(_cond_data_1538),
    .d(__muladd_madd_odata_1539)
  );

  reg [5-1:0] __delay_data_2091__delay_2090__delay_2089____variable_1522;
  reg [5-1:0] __delay_data_2092__delay_2091__delay_2090____variable_1522;
  reg [5-1:0] __delay_data_2093__delay_2092__delay_2091____variable_1522;
  reg [5-1:0] __delay_data_2094__delay_2093__delay_2092____variable_1522;
  reg signed [32-1:0] _sra_data_1540;
  wire signed [32-1:0] mul_26_z_data;
  assign mul_26_z_data = _sra_data_1540;
  wire signed [64-1:0] add_tree_16_var0_data;
  wire signed [64-1:0] add_tree_16_var1_data;
  wire signed [64-1:0] add_tree_16_var2_data;
  wire signed [64-1:0] add_tree_16_var3_data;
  wire signed [64-1:0] add_tree_16_var4_data;
  wire signed [64-1:0] add_tree_16_var5_data;
  wire signed [64-1:0] add_tree_16_var6_data;
  wire signed [64-1:0] add_tree_16_var7_data;
  wire signed [64-1:0] add_tree_16_var8_data;
  reg __add_tree_16_stream_ivalid_1;
  reg __add_tree_16_stream_ivalid_2;
  reg signed [64-1:0] __plusn_data_1314;
  reg signed [64-1:0] __plusn_data_1315;
  reg signed [64-1:0] __plusn_data_1316;
  reg signed [64-1:0] __plusn_data_1317;
  wire signed [64-1:0] add_tree_16_sum_data;
  assign add_tree_16_sum_data = __plusn_data_1317;
  wire signed [64-1:0] acc_14_x_data;
  wire [7-1:0] acc_14_rshift_data;
  wire [32-1:0] acc_14_size_data;
  wire [1-1:0] acc_14__reduce_reset_data;
  reg __acc_14_stream_ivalid_1;
  reg __acc_14_stream_ivalid_2;
  reg __acc_14_stream_ivalid_3;
  reg __acc_14_stream_ivalid_4;
  reg __acc_14_stream_ivalid_5;
  reg [1-1:0] _greaterthan_data_1283;
  reg [7-1:0] _minus_data_1285;
  reg signed [64-1:0] _reduceadd_data_1296;
  reg [33-1:0] _reduceadd_count_1296;
  reg _reduceadd_prev_count_max_1296;
  wire _reduceadd_reset_cond_1296;
  assign _reduceadd_reset_cond_1296 = acc_14__reduce_reset_data || _reduceadd_prev_count_max_1296;
  wire [33-1:0] _reduceadd_current_count_1296;
  assign _reduceadd_current_count_1296 = (_reduceadd_reset_cond_1296)? 0 : _reduceadd_count_1296;
  wire signed [64-1:0] _reduceadd_current_data_1296;
  assign _reduceadd_current_data_1296 = (_reduceadd_reset_cond_1296)? 1'sd0 : _reduceadd_data_1296;
  reg [1-1:0] _pulse_data_1298;
  reg [33-1:0] _pulse_count_1298;
  reg _pulse_prev_count_max_1298;
  wire _pulse_reset_cond_1298;
  assign _pulse_reset_cond_1298 = acc_14__reduce_reset_data || _pulse_prev_count_max_1298;
  wire [33-1:0] _pulse_current_count_1298;
  assign _pulse_current_count_1298 = (_pulse_reset_cond_1298)? 0 : _pulse_count_1298;
  wire [1-1:0] _pulse_current_data_1298;
  assign _pulse_current_data_1298 = (_pulse_reset_cond_1298)? 1'sd0 : _pulse_data_1298;
  reg [7-1:0] __delay_data_2103__variable_1281;
  reg signed [130-1:0] _sll_data_1287;
  reg [1-1:0] __delay_data_2100_greaterthan_1283;
  reg signed [64-1:0] __delay_data_2101_reduceadd_1296;
  reg [7-1:0] __delay_data_2104__delay_2103__variable_1281;
  reg [1-1:0] __delay_data_2107_pulse_1298;
  reg signed [64-1:0] _cond_data_1293;
  reg signed [64-1:0] __delay_data_2102__delay_2101_reduceadd_1296;
  reg [7-1:0] __delay_data_2105__delay_2104__delay_2103__variable_1281;
  reg [1-1:0] __delay_data_2108__delay_2107_pulse_1298;
  reg signed [64-1:0] _plus_data_1300;
  reg [7-1:0] __delay_data_2106__delay_2105__delay_2104____variable_1281;
  reg [1-1:0] __delay_data_2109__delay_2108__delay_2107_pulse_1298;
  reg signed [64-1:0] _sra_data_1301;
  reg [1-1:0] __delay_data_2110__delay_2109__delay_2108___pulse_1298;
  wire signed [64-1:0] acc_14_sum_data;
  assign acc_14_sum_data = _sra_data_1301;
  wire [1-1:0] acc_14_valid_data;
  assign acc_14_valid_data = __delay_data_2110__delay_2109__delay_2108___pulse_1298;
  wire signed [64-1:0] mul_rshift_round_clip_17_x_data;
  wire signed [16-1:0] mul_rshift_round_clip_17_y_data;
  wire [7-1:0] mul_rshift_round_clip_17_rshift_data;
  reg __mul_rshift_round_clip_17_stream_ivalid_1;
  reg __mul_rshift_round_clip_17_stream_ivalid_2;
  reg __mul_rshift_round_clip_17_stream_ivalid_3;
  reg __mul_rshift_round_clip_17_stream_ivalid_4;
  reg __mul_rshift_round_clip_17_stream_ivalid_5;
  reg __mul_rshift_round_clip_17_stream_ivalid_6;
  reg __mul_rshift_round_clip_17_stream_ivalid_7;
  reg __mul_rshift_round_clip_17_stream_ivalid_8;
  wire signed [80-1:0] _times_mul_odata_1321;
  reg signed [80-1:0] _times_mul_odata_reg_1321;
  wire signed [80-1:0] _times_data_1321;
  assign _times_data_1321 = _times_mul_odata_reg_1321;
  wire _times_mul_update_1321;
  assign _times_mul_update_1321 = _mul_rshift_round_clip_17_stream_oready;

  multiplier_1
  _times_mul_1321
  (
    .CLK(CLK),
    .update(_times_mul_update_1321),
    .a(mul_rshift_round_clip_17_x_data),
    .b(mul_rshift_round_clip_17_y_data),
    .c(_times_mul_odata_1321)
  );

  wire [7-1:0] _minus_data_1324;
  assign _minus_data_1324 = mul_rshift_round_clip_17_rshift_data - 2'sd1;
  wire signed [130-1:0] _sll_data_1327;
  assign _sll_data_1327 = 2'sd1 << _minus_data_1324;
  wire [1-1:0] _eq_data_1339;
  assign _eq_data_1339 = mul_rshift_round_clip_17_rshift_data == 1'sd0;
  reg signed [130-1:0] __delay_data_2116_sll_1327;
  reg [7-1:0] __delay_data_2120__variable_1320;
  reg [1-1:0] __delay_data_2124_eq_1339;
  reg signed [130-1:0] __delay_data_2117__delay_2116_sll_1327;
  reg [7-1:0] __delay_data_2121__delay_2120__variable_1320;
  reg [1-1:0] __delay_data_2125__delay_2124_eq_1339;
  reg signed [130-1:0] __delay_data_2118__delay_2117__delay_2116_sll_1327;
  reg [7-1:0] __delay_data_2122__delay_2121__delay_2120__variable_1320;
  reg [1-1:0] __delay_data_2126__delay_2125__delay_2124_eq_1339;
  reg signed [130-1:0] __delay_data_2119__delay_2118__delay_2117__delay_2116_sll_1327;
  reg [7-1:0] __delay_data_2123__delay_2122__delay_2121____variable_1320;
  reg [1-1:0] __delay_data_2127__delay_2126__delay_2125__delay_2124_eq_1339;
  wire [1-1:0] _pointer_data_1322;
  assign _pointer_data_1322 = _times_data_1321[8'sd79];
  wire signed [2-1:0] _cond_data_1334;
  assign _cond_data_1334 = (_pointer_data_1322)? -2'sd1 : 1'sd0;
  wire signed [81-1:0] _plus_data_1335;
  assign _plus_data_1335 = _times_data_1321 + __delay_data_2119__delay_2118__delay_2117__delay_2116_sll_1327;
  wire signed [81-1:0] _plus_data_1336;
  assign _plus_data_1336 = _plus_data_1335 + _cond_data_1334;
  wire signed [80-1:0] _sra_data_1337;
  assign _sra_data_1337 = _plus_data_1336 >>> __delay_data_2123__delay_2122__delay_2121____variable_1320;
  reg signed [80-1:0] _cond_data_1340;
  reg [1-1:0] _greaterthan_data_1341;
  reg [1-1:0] _lessthan_data_1345;
  reg [1-1:0] _greatereq_data_1349;
  reg signed [80-1:0] __delay_data_2128_cond_1340;
  reg signed [80-1:0] _cond_data_1343;
  reg signed [80-1:0] _cond_data_1347;
  reg [1-1:0] __delay_data_2129_greatereq_1349;
  reg signed [16-1:0] _cond_data_1351;
  wire signed [16-1:0] mul_rshift_round_clip_17_z_data;
  assign mul_rshift_round_clip_17_z_data = _cond_data_1351;
  reg [33-1:0] _stream_conv2d_4_sink_50_sink_count;
  reg [5-1:0] _stream_conv2d_4_sink_50_sink_mode;
  reg [16-1:0] _stream_conv2d_4_sink_50_sink_generator_id;
  reg [32-1:0] _stream_conv2d_4_sink_50_sink_offset;
  reg [33-1:0] _stream_conv2d_4_sink_50_sink_size;
  reg [32-1:0] _stream_conv2d_4_sink_50_sink_stride;
  reg [32-1:0] _stream_conv2d_4_sink_50_sink_offset_buf;
  reg [33-1:0] _stream_conv2d_4_sink_50_sink_size_buf;
  reg [32-1:0] _stream_conv2d_4_sink_50_sink_stride_buf;
  reg [8-1:0] _stream_conv2d_4_sink_50_sink_sel;
  reg [32-1:0] _stream_conv2d_4_sink_50_sink_waddr;
  reg _stream_conv2d_4_sink_50_sink_wenable;
  reg [16-1:0] _stream_conv2d_4_sink_50_sink_wdata;
  reg _stream_conv2d_4_sink_50_sink_fifo_enq;
  reg [16-1:0] _stream_conv2d_4_sink_50_sink_fifo_wdata;
  reg [16-1:0] _stream_conv2d_4_sink_50_sink_immediate;
  reg [33-1:0] _stream_conv2d_4_sink_51_sink_count;
  reg [5-1:0] _stream_conv2d_4_sink_51_sink_mode;
  reg [16-1:0] _stream_conv2d_4_sink_51_sink_generator_id;
  reg [32-1:0] _stream_conv2d_4_sink_51_sink_offset;
  reg [33-1:0] _stream_conv2d_4_sink_51_sink_size;
  reg [32-1:0] _stream_conv2d_4_sink_51_sink_stride;
  reg [32-1:0] _stream_conv2d_4_sink_51_sink_offset_buf;
  reg [33-1:0] _stream_conv2d_4_sink_51_sink_size_buf;
  reg [32-1:0] _stream_conv2d_4_sink_51_sink_stride_buf;
  reg [8-1:0] _stream_conv2d_4_sink_51_sink_sel;
  reg [32-1:0] _stream_conv2d_4_sink_51_sink_waddr;
  reg _stream_conv2d_4_sink_51_sink_wenable;
  reg [1-1:0] _stream_conv2d_4_sink_51_sink_wdata;
  reg _stream_conv2d_4_sink_51_sink_fifo_enq;
  reg [1-1:0] _stream_conv2d_4_sink_51_sink_fifo_wdata;
  reg [1-1:0] _stream_conv2d_4_sink_51_sink_immediate;
  reg _stream_max_pool_serial_6_stream_ivalid;
  wire _stream_max_pool_serial_6_stream_oready;
  wire _stream_max_pool_serial_6_stream_internal_oready;
  assign _stream_max_pool_serial_6_stream_oready = _stream_max_pool_serial_6_stream_internal_oready;
  reg [32-1:0] _stream_max_pool_serial_6_fsm;
  localparam _stream_max_pool_serial_6_fsm_init = 0;
  wire _stream_max_pool_serial_6_run_flag;
  reg _stream_max_pool_serial_6_source_start;
  wire _stream_max_pool_serial_6_source_stop;
  reg _stream_max_pool_serial_6_source_busy;
  wire _stream_max_pool_serial_6_sink_start;
  wire _stream_max_pool_serial_6_sink_stop;
  wire _stream_max_pool_serial_6_sink_busy;
  wire _stream_max_pool_serial_6_busy;
  reg _stream_max_pool_serial_6_busy_reg;
  wire _stream_max_pool_serial_6_is_root;
  assign _stream_max_pool_serial_6_is_root = 1;
  reg [3-1:0] _stream_max_pool_serial_6_parameter_0_next_parameter_data;
  reg _stream_max_pool_serial_6_source_1_idle;
  reg [33-1:0] _stream_max_pool_serial_6_source_1_source_count;
  reg [5-1:0] _stream_max_pool_serial_6_source_1_source_mode;
  reg [16-1:0] _stream_max_pool_serial_6_source_1_source_generator_id;
  reg [32-1:0] _stream_max_pool_serial_6_source_1_source_offset;
  reg [33-1:0] _stream_max_pool_serial_6_source_1_source_size;
  reg [32-1:0] _stream_max_pool_serial_6_source_1_source_stride;
  reg [32-1:0] _stream_max_pool_serial_6_source_1_source_offset_buf;
  reg [33-1:0] _stream_max_pool_serial_6_source_1_source_size_buf;
  reg [32-1:0] _stream_max_pool_serial_6_source_1_source_stride_buf;
  reg [8-1:0] _stream_max_pool_serial_6_source_1_source_sel;
  reg [32-1:0] _stream_max_pool_serial_6_source_1_source_ram_raddr;
  reg _stream_max_pool_serial_6_source_1_source_ram_renable;
  wire [16-1:0] _stream_max_pool_serial_6_source_1_source_ram_rdata;
  reg _stream_max_pool_serial_6_source_1_source_fifo_deq;
  wire [16-1:0] _stream_max_pool_serial_6_source_1_source_fifo_rdata;
  reg [16-1:0] _stream_max_pool_serial_6_source_1_source_empty_data;
  reg [4-1:0] _stream_max_pool_serial_6_parameter_2_next_parameter_data;
  wire signed [16-1:0] _reduce_max_27_x_data;
  wire [32-1:0] _reduce_max_27_size_data;
  wire [1-1:0] _reduce_max_27__reduce_reset_data;
  reg ___reduce_max_27_stream_ivalid_1;
  reg signed [16-1:0] _reducemax_data_1544;
  reg [33-1:0] _reducemax_count_1544;
  reg _reducemax_prev_count_max_1544;
  wire _reducemax_reset_cond_1544;
  assign _reducemax_reset_cond_1544 = _reduce_max_27__reduce_reset_data || _reducemax_prev_count_max_1544;
  wire [33-1:0] _reducemax_current_count_1544;
  assign _reducemax_current_count_1544 = (_reducemax_reset_cond_1544)? 0 : _reducemax_count_1544;
  wire signed [16-1:0] _reducemax_current_data_1544;
  assign _reducemax_current_data_1544 = (_reducemax_reset_cond_1544)? -17'sd32768 : _reducemax_data_1544;
  reg [1-1:0] _pulse_data_1546;
  reg [33-1:0] _pulse_count_1546;
  reg _pulse_prev_count_max_1546;
  wire _pulse_reset_cond_1546;
  assign _pulse_reset_cond_1546 = _reduce_max_27__reduce_reset_data || _pulse_prev_count_max_1546;
  wire [33-1:0] _pulse_current_count_1546;
  assign _pulse_current_count_1546 = (_pulse_reset_cond_1546)? 0 : _pulse_count_1546;
  wire [1-1:0] _pulse_current_data_1546;
  assign _pulse_current_data_1546 = (_pulse_reset_cond_1546)? 1'sd0 : _pulse_data_1546;
  wire signed [16-1:0] _reduce_max_27_data_data;
  assign _reduce_max_27_data_data = _reducemax_data_1544;
  wire [1-1:0] _reduce_max_27_valid_data;
  assign _reduce_max_27_valid_data = _pulse_data_1546;
  reg [33-1:0] _stream_max_pool_serial_6_sink_5_sink_count;
  reg [5-1:0] _stream_max_pool_serial_6_sink_5_sink_mode;
  reg [16-1:0] _stream_max_pool_serial_6_sink_5_sink_generator_id;
  reg [32-1:0] _stream_max_pool_serial_6_sink_5_sink_offset;
  reg [33-1:0] _stream_max_pool_serial_6_sink_5_sink_size;
  reg [32-1:0] _stream_max_pool_serial_6_sink_5_sink_stride;
  reg [32-1:0] _stream_max_pool_serial_6_sink_5_sink_offset_buf;
  reg [33-1:0] _stream_max_pool_serial_6_sink_5_sink_size_buf;
  reg [32-1:0] _stream_max_pool_serial_6_sink_5_sink_stride_buf;
  reg [8-1:0] _stream_max_pool_serial_6_sink_5_sink_sel;
  reg [32-1:0] _stream_max_pool_serial_6_sink_5_sink_waddr;
  reg _stream_max_pool_serial_6_sink_5_sink_wenable;
  reg [16-1:0] _stream_max_pool_serial_6_sink_5_sink_wdata;
  reg _stream_max_pool_serial_6_sink_5_sink_fifo_enq;
  reg [16-1:0] _stream_max_pool_serial_6_sink_5_sink_fifo_wdata;
  reg [16-1:0] _stream_max_pool_serial_6_sink_5_sink_immediate;
  reg [33-1:0] _stream_max_pool_serial_6_sink_6_sink_count;
  reg [5-1:0] _stream_max_pool_serial_6_sink_6_sink_mode;
  reg [16-1:0] _stream_max_pool_serial_6_sink_6_sink_generator_id;
  reg [32-1:0] _stream_max_pool_serial_6_sink_6_sink_offset;
  reg [33-1:0] _stream_max_pool_serial_6_sink_6_sink_size;
  reg [32-1:0] _stream_max_pool_serial_6_sink_6_sink_stride;
  reg [32-1:0] _stream_max_pool_serial_6_sink_6_sink_offset_buf;
  reg [33-1:0] _stream_max_pool_serial_6_sink_6_sink_size_buf;
  reg [32-1:0] _stream_max_pool_serial_6_sink_6_sink_stride_buf;
  reg [8-1:0] _stream_max_pool_serial_6_sink_6_sink_sel;
  reg [32-1:0] _stream_max_pool_serial_6_sink_6_sink_waddr;
  reg _stream_max_pool_serial_6_sink_6_sink_wenable;
  reg [1-1:0] _stream_max_pool_serial_6_sink_6_sink_wdata;
  reg _stream_max_pool_serial_6_sink_6_sink_fifo_enq;
  reg [1-1:0] _stream_max_pool_serial_6_sink_6_sink_fifo_wdata;
  reg [1-1:0] _stream_max_pool_serial_6_sink_6_sink_immediate;
  reg _stream_matmul_11_stream_ivalid;
  wire _stream_matmul_11_stream_oready;
  wire _stream_matmul_11_stream_internal_oready;
  assign _stream_matmul_11_stream_oready = _stream_matmul_11_stream_internal_oready;
  reg [32-1:0] _stream_matmul_11_fsm;
  localparam _stream_matmul_11_fsm_init = 0;
  wire _stream_matmul_11_run_flag;
  reg _stream_matmul_11_source_start;
  wire _stream_matmul_11_source_stop;
  reg _stream_matmul_11_source_busy;
  wire _stream_matmul_11_sink_start;
  wire _stream_matmul_11_sink_stop;
  wire _stream_matmul_11_sink_busy;
  wire _stream_matmul_11_busy;
  reg _stream_matmul_11_busy_reg;
  wire _stream_matmul_11_is_root;
  assign _stream_matmul_11_is_root = 1;
  reg [13-1:0] _stream_matmul_11_parameter_0_next_parameter_data;
  reg [1-1:0] _stream_matmul_11_parameter_1_next_parameter_data;
  reg [1-1:0] _stream_matmul_11_parameter_2_next_parameter_data;
  reg [1-1:0] _stream_matmul_11_parameter_3_next_parameter_data;
  reg [1-1:0] _stream_matmul_11_parameter_4_next_parameter_data;
  reg [1-1:0] _stream_matmul_11_parameter_6_next_parameter_data;
  reg _stream_matmul_11_source_7_idle;
  reg [33-1:0] _stream_matmul_11_source_7_source_count;
  reg [5-1:0] _stream_matmul_11_source_7_source_mode;
  reg [16-1:0] _stream_matmul_11_source_7_source_generator_id;
  reg [32-1:0] _stream_matmul_11_source_7_source_offset;
  reg [33-1:0] _stream_matmul_11_source_7_source_size;
  reg [32-1:0] _stream_matmul_11_source_7_source_stride;
  reg [32-1:0] _stream_matmul_11_source_7_source_offset_buf;
  reg [33-1:0] _stream_matmul_11_source_7_source_size_buf;
  reg [32-1:0] _stream_matmul_11_source_7_source_stride_buf;
  reg [8-1:0] _stream_matmul_11_source_7_source_sel;
  reg [32-1:0] _stream_matmul_11_source_7_source_ram_raddr;
  reg _stream_matmul_11_source_7_source_ram_renable;
  wire [16-1:0] _stream_matmul_11_source_7_source_ram_rdata;
  reg _stream_matmul_11_source_7_source_fifo_deq;
  wire [16-1:0] _stream_matmul_11_source_7_source_fifo_rdata;
  reg [16-1:0] _stream_matmul_11_source_7_source_empty_data;
  reg [1-1:0] _stream_matmul_11_parameter_8_next_parameter_data;
  reg _stream_matmul_11_source_9_idle;
  reg [33-1:0] _stream_matmul_11_source_9_source_count;
  reg [5-1:0] _stream_matmul_11_source_9_source_mode;
  reg [16-1:0] _stream_matmul_11_source_9_source_generator_id;
  reg [32-1:0] _stream_matmul_11_source_9_source_offset;
  reg [33-1:0] _stream_matmul_11_source_9_source_size;
  reg [32-1:0] _stream_matmul_11_source_9_source_stride;
  reg [32-1:0] _stream_matmul_11_source_9_source_offset_buf;
  reg [33-1:0] _stream_matmul_11_source_9_source_size_buf;
  reg [32-1:0] _stream_matmul_11_source_9_source_stride_buf;
  reg [8-1:0] _stream_matmul_11_source_9_source_sel;
  reg [32-1:0] _stream_matmul_11_source_9_source_ram_raddr;
  reg _stream_matmul_11_source_9_source_ram_renable;
  wire [16-1:0] _stream_matmul_11_source_9_source_ram_rdata;
  reg _stream_matmul_11_source_9_source_fifo_deq;
  wire [16-1:0] _stream_matmul_11_source_9_source_fifo_rdata;
  reg [16-1:0] _stream_matmul_11_source_9_source_empty_data;
  reg [1-1:0] _stream_matmul_11_parameter_10_next_parameter_data;
  reg _stream_matmul_11_source_11_idle;
  reg [33-1:0] _stream_matmul_11_source_11_source_count;
  reg [5-1:0] _stream_matmul_11_source_11_source_mode;
  reg [16-1:0] _stream_matmul_11_source_11_source_generator_id;
  reg [32-1:0] _stream_matmul_11_source_11_source_offset;
  reg [33-1:0] _stream_matmul_11_source_11_source_size;
  reg [32-1:0] _stream_matmul_11_source_11_source_stride;
  reg [32-1:0] _stream_matmul_11_source_11_source_offset_buf;
  reg [33-1:0] _stream_matmul_11_source_11_source_size_buf;
  reg [32-1:0] _stream_matmul_11_source_11_source_stride_buf;
  reg [8-1:0] _stream_matmul_11_source_11_source_sel;
  reg [32-1:0] _stream_matmul_11_source_11_source_ram_raddr;
  reg _stream_matmul_11_source_11_source_ram_renable;
  wire [16-1:0] _stream_matmul_11_source_11_source_ram_rdata;
  reg _stream_matmul_11_source_11_source_fifo_deq;
  wire [16-1:0] _stream_matmul_11_source_11_source_fifo_rdata;
  reg [16-1:0] _stream_matmul_11_source_11_source_empty_data;
  reg [1-1:0] _stream_matmul_11_parameter_12_next_parameter_data;
  reg _stream_matmul_11_source_13_idle;
  reg [33-1:0] _stream_matmul_11_source_13_source_count;
  reg [5-1:0] _stream_matmul_11_source_13_source_mode;
  reg [16-1:0] _stream_matmul_11_source_13_source_generator_id;
  reg [32-1:0] _stream_matmul_11_source_13_source_offset;
  reg [33-1:0] _stream_matmul_11_source_13_source_size;
  reg [32-1:0] _stream_matmul_11_source_13_source_stride;
  reg [32-1:0] _stream_matmul_11_source_13_source_offset_buf;
  reg [33-1:0] _stream_matmul_11_source_13_source_size_buf;
  reg [32-1:0] _stream_matmul_11_source_13_source_stride_buf;
  reg [8-1:0] _stream_matmul_11_source_13_source_sel;
  reg [32-1:0] _stream_matmul_11_source_13_source_ram_raddr;
  reg _stream_matmul_11_source_13_source_ram_renable;
  wire [16-1:0] _stream_matmul_11_source_13_source_ram_rdata;
  reg _stream_matmul_11_source_13_source_fifo_deq;
  wire [16-1:0] _stream_matmul_11_source_13_source_fifo_rdata;
  reg [16-1:0] _stream_matmul_11_source_13_source_empty_data;
  reg [1-1:0] _stream_matmul_11_parameter_14_next_parameter_data;
  reg _stream_matmul_11_source_15_idle;
  reg [33-1:0] _stream_matmul_11_source_15_source_count;
  reg [5-1:0] _stream_matmul_11_source_15_source_mode;
  reg [16-1:0] _stream_matmul_11_source_15_source_generator_id;
  reg [32-1:0] _stream_matmul_11_source_15_source_offset;
  reg [33-1:0] _stream_matmul_11_source_15_source_size;
  reg [32-1:0] _stream_matmul_11_source_15_source_stride;
  reg [32-1:0] _stream_matmul_11_source_15_source_offset_buf;
  reg [33-1:0] _stream_matmul_11_source_15_source_size_buf;
  reg [32-1:0] _stream_matmul_11_source_15_source_stride_buf;
  reg [8-1:0] _stream_matmul_11_source_15_source_sel;
  reg [32-1:0] _stream_matmul_11_source_15_source_ram_raddr;
  reg _stream_matmul_11_source_15_source_ram_renable;
  wire [16-1:0] _stream_matmul_11_source_15_source_ram_rdata;
  reg _stream_matmul_11_source_15_source_fifo_deq;
  wire [16-1:0] _stream_matmul_11_source_15_source_fifo_rdata;
  reg [16-1:0] _stream_matmul_11_source_15_source_empty_data;
  reg [1-1:0] _stream_matmul_11_parameter_16_next_parameter_data;
  reg [1-1:0] _stream_matmul_11_parameter_17_next_parameter_data;
  reg [5-1:0] _stream_matmul_11_parameter_18_next_parameter_data;
  reg [2-1:0] _stream_matmul_11_parameter_19_next_parameter_data;
  reg _stream_matmul_11_source_20_idle;
  reg [33-1:0] _stream_matmul_11_source_20_source_count;
  reg [5-1:0] _stream_matmul_11_source_20_source_mode;
  reg [16-1:0] _stream_matmul_11_source_20_source_generator_id;
  reg [32-1:0] _stream_matmul_11_source_20_source_offset;
  reg [33-1:0] _stream_matmul_11_source_20_source_size;
  reg [32-1:0] _stream_matmul_11_source_20_source_stride;
  reg [32-1:0] _stream_matmul_11_source_20_source_offset_buf;
  reg [33-1:0] _stream_matmul_11_source_20_source_size_buf;
  reg [32-1:0] _stream_matmul_11_source_20_source_stride_buf;
  reg [8-1:0] _stream_matmul_11_source_20_source_sel;
  reg [32-1:0] _stream_matmul_11_source_20_source_ram_raddr;
  reg _stream_matmul_11_source_20_source_ram_renable;
  wire [16-1:0] _stream_matmul_11_source_20_source_ram_rdata;
  reg _stream_matmul_11_source_20_source_fifo_deq;
  wire [16-1:0] _stream_matmul_11_source_20_source_fifo_rdata;
  reg [16-1:0] _stream_matmul_11_source_20_source_empty_data;
  reg _stream_matmul_11_source_21_idle;
  reg [33-1:0] _stream_matmul_11_source_21_source_count;
  reg [5-1:0] _stream_matmul_11_source_21_source_mode;
  reg [16-1:0] _stream_matmul_11_source_21_source_generator_id;
  reg [32-1:0] _stream_matmul_11_source_21_source_offset;
  reg [33-1:0] _stream_matmul_11_source_21_source_size;
  reg [32-1:0] _stream_matmul_11_source_21_source_stride;
  reg [32-1:0] _stream_matmul_11_source_21_source_offset_buf;
  reg [33-1:0] _stream_matmul_11_source_21_source_size_buf;
  reg [32-1:0] _stream_matmul_11_source_21_source_stride_buf;
  reg [8-1:0] _stream_matmul_11_source_21_source_sel;
  reg [32-1:0] _stream_matmul_11_source_21_source_ram_raddr;
  reg _stream_matmul_11_source_21_source_ram_renable;
  wire [16-1:0] _stream_matmul_11_source_21_source_ram_rdata;
  reg _stream_matmul_11_source_21_source_fifo_deq;
  wire [16-1:0] _stream_matmul_11_source_21_source_fifo_rdata;
  reg [16-1:0] _stream_matmul_11_source_21_source_empty_data;
  wire signed [64-1:0] add_tree_15_var0_data;
  wire signed [64-1:0] _cast_src_1303;
  assign _cast_src_1303 = add_tree_15_var0_data;
  wire signed [64-1:0] _cast_data_1303;
  assign _cast_data_1303 = _cast_src_1303;
  wire signed [64-1:0] add_tree_15_sum_data;
  assign add_tree_15_sum_data = _cast_data_1303;
  reg [33-1:0] _stream_matmul_11_sink_26_sink_count;
  reg [5-1:0] _stream_matmul_11_sink_26_sink_mode;
  reg [16-1:0] _stream_matmul_11_sink_26_sink_generator_id;
  reg [32-1:0] _stream_matmul_11_sink_26_sink_offset;
  reg [33-1:0] _stream_matmul_11_sink_26_sink_size;
  reg [32-1:0] _stream_matmul_11_sink_26_sink_stride;
  reg [32-1:0] _stream_matmul_11_sink_26_sink_offset_buf;
  reg [33-1:0] _stream_matmul_11_sink_26_sink_size_buf;
  reg [32-1:0] _stream_matmul_11_sink_26_sink_stride_buf;
  reg [8-1:0] _stream_matmul_11_sink_26_sink_sel;
  reg [32-1:0] _stream_matmul_11_sink_26_sink_waddr;
  reg _stream_matmul_11_sink_26_sink_wenable;
  reg [16-1:0] _stream_matmul_11_sink_26_sink_wdata;
  reg _stream_matmul_11_sink_26_sink_fifo_enq;
  reg [16-1:0] _stream_matmul_11_sink_26_sink_fifo_wdata;
  reg [16-1:0] _stream_matmul_11_sink_26_sink_immediate;
  reg [33-1:0] _stream_matmul_11_sink_27_sink_count;
  reg [5-1:0] _stream_matmul_11_sink_27_sink_mode;
  reg [16-1:0] _stream_matmul_11_sink_27_sink_generator_id;
  reg [32-1:0] _stream_matmul_11_sink_27_sink_offset;
  reg [33-1:0] _stream_matmul_11_sink_27_sink_size;
  reg [32-1:0] _stream_matmul_11_sink_27_sink_stride;
  reg [32-1:0] _stream_matmul_11_sink_27_sink_offset_buf;
  reg [33-1:0] _stream_matmul_11_sink_27_sink_size_buf;
  reg [32-1:0] _stream_matmul_11_sink_27_sink_stride_buf;
  reg [8-1:0] _stream_matmul_11_sink_27_sink_sel;
  reg [32-1:0] _stream_matmul_11_sink_27_sink_waddr;
  reg _stream_matmul_11_sink_27_sink_wenable;
  reg [1-1:0] _stream_matmul_11_sink_27_sink_wdata;
  reg _stream_matmul_11_sink_27_sink_fifo_enq;
  reg [1-1:0] _stream_matmul_11_sink_27_sink_fifo_wdata;
  reg [1-1:0] _stream_matmul_11_sink_27_sink_immediate;
  reg [32-1:0] main_fsm;
  localparam main_fsm_init = 0;
  reg [32-1:0] internal_state_counter;
  reg [32-1:0] conv2d_4_objaddr;
  reg [32-1:0] conv2d_4_arg_objaddr_0;
  reg [32-1:0] conv2d_4_arg_objaddr_1;
  reg [32-1:0] conv2d_4_arg_objaddr_2;
  reg [32-1:0] conv2d_4_arg_objaddr_3;
  reg [32-1:0] control_conv2d_4;
  localparam control_conv2d_4_init = 0;
  reg _control_conv2d_4_called;
  wire signed [32-1:0] conv2d_4_act_base_offset;
  reg signed [32-1:0] conv2d_4_act_base_offset_row;
  reg signed [32-1:0] conv2d_4_act_base_offset_bat;
  assign conv2d_4_act_base_offset = conv2d_4_act_base_offset_row + conv2d_4_act_base_offset_bat;
  reg signed [32-1:0] conv2d_4_filter_base_offset;
  reg [32-1:0] conv2d_4_next_stream_num_ops;
  wire signed [32-1:0] conv2d_4_out_base_offset;
  reg signed [32-1:0] conv2d_4_out_base_offset_val;
  reg signed [32-1:0] conv2d_4_out_base_offset_col;
  reg signed [32-1:0] conv2d_4_out_base_offset_row;
  reg signed [32-1:0] conv2d_4_out_base_offset_bat;
  reg signed [32-1:0] conv2d_4_out_base_offset_och;
  assign conv2d_4_out_base_offset = conv2d_4_out_base_offset_val + conv2d_4_out_base_offset_col + conv2d_4_out_base_offset_row + conv2d_4_out_base_offset_bat + conv2d_4_out_base_offset_och;
  reg conv2d_4_dma_flag_0;
  reg conv2d_4_dma_flag_1;
  reg conv2d_4_dma_flag_2;
  reg [32-1:0] conv2d_4_sync_comp_count;
  reg [32-1:0] conv2d_4_sync_out_count;
  reg [32-1:0] conv2d_4_write_count;
  reg [32-1:0] conv2d_4_next_out_write_size;
  reg [32-1:0] conv2d_4_col_count;
  reg [32-1:0] conv2d_4_row_count;
  reg [32-1:0] conv2d_4_bat_count;
  reg [32-1:0] conv2d_4_och_count;
  reg [2-1:0] conv2d_4_col_select;
  reg [2-1:0] conv2d_4_row_select;
  reg [32-1:0] conv2d_4_out_col_count;
  reg [32-1:0] conv2d_4_out_row_count;
  reg [32-1:0] conv2d_4_out_ram_select;
  reg [32-1:0] conv2d_4_prev_col_count;
  reg [32-1:0] conv2d_4_prev_row_count;
  reg [32-1:0] conv2d_4_prev_bat_count;
  reg [32-1:0] conv2d_4_prev_och_count;
  reg [2-1:0] conv2d_4_prev_row_select;
  reg [32-1:0] conv2d_4_stream_act_local_0;
  reg [32-1:0] conv2d_4_stream_act_local_1;
  reg [32-1:0] conv2d_4_stream_act_local_2;
  reg [32-1:0] conv2d_4_stream_act_local_3;
  reg [32-1:0] conv2d_4_stream_act_local_4;
  reg [32-1:0] conv2d_4_stream_act_local_5;
  reg [32-1:0] conv2d_4_stream_act_local_6;
  reg [32-1:0] conv2d_4_stream_act_local_7;
  reg [32-1:0] conv2d_4_stream_act_local_8;
  reg [32-1:0] conv2d_4_stream_out_local_val;
  reg [32-1:0] conv2d_4_stream_out_local_col;
  wire [32-1:0] conv2d_4_stream_out_local;
  assign conv2d_4_stream_out_local = conv2d_4_stream_out_local_val + conv2d_4_stream_out_local_col;
  reg [32-1:0] conv2d_4_act_page_comp_offset_0;
  reg [32-1:0] conv2d_4_act_page_comp_offset_1;
  reg [32-1:0] conv2d_4_act_page_comp_offset_2;
  reg [32-1:0] conv2d_4_act_page_dma_offset_0;
  reg [32-1:0] conv2d_4_act_page_dma_offset_1;
  reg [32-1:0] conv2d_4_act_page_dma_offset_2;
  reg [32-1:0] conv2d_4_filter_page_comp_offset;
  reg [32-1:0] conv2d_4_filter_page_dma_offset;
  reg conv2d_4_out_page;
  reg [32-1:0] conv2d_4_out_page_comp_offset;
  reg [32-1:0] conv2d_4_out_page_dma_offset;
  reg [32-1:0] conv2d_4_out_laddr_offset;
  reg conv2d_4_skip_read_filter;
  reg conv2d_4_skip_read_act;
  reg conv2d_4_skip_comp;
  reg conv2d_4_skip_write_out;
  wire [6-1:0] _dma_read_packed_high_local_size_54;
  assign _dma_read_packed_high_local_size_54 = cparam_conv2d_4_bias_num >> 1;
  wire [1-1:0] _dma_read_packed_low_local_size_55;
  assign _dma_read_packed_low_local_size_55 = cparam_conv2d_4_bias_num & { 1{ 1'd1 } };
  wire [6-1:0] _dma_read_packed_local_packed_size_56;
  assign _dma_read_packed_local_packed_size_56 = (_dma_read_packed_low_local_size_55 > 0)? _dma_read_packed_high_local_size_54 + 1 : _dma_read_packed_high_local_size_54;
  wire [32-1:0] mask_addr_shifted_57;
  assign mask_addr_shifted_57 = conv2d_4_arg_objaddr_2 + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_58;
  assign mask_addr_masked_58 = mask_addr_shifted_57 << 2;
  reg [32-1:0] _maxi_read_req_fsm;
  localparam _maxi_read_req_fsm_init = 0;
  reg [33-1:0] _maxi_read_cur_global_size;
  reg _maxi_read_cont;
  wire [8-1:0] pack_read_req_op_sel_59;
  wire [32-1:0] pack_read_req_local_addr_60;
  wire [32-1:0] pack_read_req_local_stride_61;
  wire [33-1:0] pack_read_req_local_size_62;
  wire [32-1:0] pack_read_req_local_blocksize_63;
  assign pack_read_req_op_sel_59 = _maxi_read_op_sel;
  assign pack_read_req_local_addr_60 = _maxi_read_local_addr;
  assign pack_read_req_local_stride_61 = _maxi_read_local_stride;
  assign pack_read_req_local_size_62 = _maxi_read_local_size;
  assign pack_read_req_local_blocksize_63 = _maxi_read_local_blocksize;
  wire [137-1:0] pack_read_req_packed_64;
  assign pack_read_req_packed_64 = { pack_read_req_op_sel_59, pack_read_req_local_addr_60, pack_read_req_local_stride_61, pack_read_req_local_size_62, pack_read_req_local_blocksize_63 };
  assign _maxi_read_req_fifo_wdata = ((_maxi_read_req_fsm == 0) && _maxi_read_start && !_maxi_read_req_fifo_almost_full)? pack_read_req_packed_64 : 'hx;
  assign _maxi_read_req_fifo_enq = ((_maxi_read_req_fsm == 0) && _maxi_read_start && !_maxi_read_req_fifo_almost_full)? (_maxi_read_req_fsm == 0) && _maxi_read_start && !_maxi_read_req_fifo_almost_full && !_maxi_read_req_fifo_almost_full : 0;
  localparam _tmp_65 = 1;
  wire [_tmp_65-1:0] _tmp_66;
  assign _tmp_66 = !_maxi_read_req_fifo_almost_full;
  reg [_tmp_65-1:0] __tmp_66_1;
  wire [32-1:0] mask_addr_shifted_67;
  assign mask_addr_shifted_67 = _maxi_read_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_68;
  assign mask_addr_masked_68 = mask_addr_shifted_67 << 2;
  wire [32-1:0] mask_addr_shifted_69;
  assign mask_addr_shifted_69 = _maxi_read_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_70;
  assign mask_addr_masked_70 = mask_addr_shifted_69 << 2;
  wire [32-1:0] mask_addr_shifted_71;
  assign mask_addr_shifted_71 = _maxi_read_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_72;
  assign mask_addr_masked_72 = mask_addr_shifted_71 << 2;
  wire [32-1:0] mask_addr_shifted_73;
  assign mask_addr_shifted_73 = _maxi_read_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_74;
  assign mask_addr_masked_74 = mask_addr_shifted_73 << 2;
  wire [32-1:0] mask_addr_shifted_75;
  assign mask_addr_shifted_75 = _maxi_read_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_76;
  assign mask_addr_masked_76 = mask_addr_shifted_75 << 2;
  wire [32-1:0] mask_addr_shifted_77;
  assign mask_addr_shifted_77 = _maxi_read_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_78;
  assign mask_addr_masked_78 = mask_addr_shifted_77 << 2;
  reg _maxi_raddr_cond_0_1;
  reg [32-1:0] _maxi_read_data_fsm;
  localparam _maxi_read_data_fsm_init = 0;
  reg [32-1:0] write_burst_packed_fsm_31;
  localparam write_burst_packed_fsm_31_init = 0;
  reg [9-1:0] write_burst_packed_addr_79;
  reg [9-1:0] write_burst_packed_stride_80;
  reg [33-1:0] write_burst_packed_length_81;
  reg write_burst_packed_done_82;
  wire [8-1:0] write_burst_packed_ram_addr_83;
  assign write_burst_packed_ram_addr_83 = write_burst_packed_addr_79 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_84;
  assign write_burst_packed_ram_wdata_84 = _maxi_rdata_sb_0 >> 0;
  assign ram_w16_l512_id9_0_1_addr = ((write_burst_packed_fsm_31 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_addr_83 : 'hx;
  assign ram_w16_l512_id9_0_1_wdata = ((write_burst_packed_fsm_31 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_wdata_84 : 'hx;
  assign ram_w16_l512_id9_0_1_wenable = ((write_burst_packed_fsm_31 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  assign ram_w16_l512_id9_0_1_enable = ((write_burst_packed_fsm_31 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  wire [8-1:0] write_burst_packed_ram_addr_85;
  assign write_burst_packed_ram_addr_85 = write_burst_packed_addr_79 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_86;
  assign write_burst_packed_ram_wdata_86 = _maxi_rdata_sb_0 >> 16;
  assign ram_w16_l512_id9_1_1_addr = ((write_burst_packed_fsm_31 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_addr_85 : 'hx;
  assign ram_w16_l512_id9_1_1_wdata = ((write_burst_packed_fsm_31 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_wdata_86 : 'hx;
  assign ram_w16_l512_id9_1_1_wenable = ((write_burst_packed_fsm_31 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  assign ram_w16_l512_id9_1_1_enable = ((write_burst_packed_fsm_31 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  wire [6-1:0] _dma_read_packed_high_local_size_87;
  assign _dma_read_packed_high_local_size_87 = cparam_conv2d_4_scale_num >> 1;
  wire [1-1:0] _dma_read_packed_low_local_size_88;
  assign _dma_read_packed_low_local_size_88 = cparam_conv2d_4_scale_num & { 1{ 1'd1 } };
  wire [6-1:0] _dma_read_packed_local_packed_size_89;
  assign _dma_read_packed_local_packed_size_89 = (_dma_read_packed_low_local_size_88 > 0)? _dma_read_packed_high_local_size_87 + 1 : _dma_read_packed_high_local_size_87;
  wire [32-1:0] mask_addr_shifted_90;
  assign mask_addr_shifted_90 = conv2d_4_arg_objaddr_3 + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_91;
  assign mask_addr_masked_91 = mask_addr_shifted_90 << 2;
  reg [32-1:0] write_burst_packed_fsm_32;
  localparam write_burst_packed_fsm_32_init = 0;
  reg [9-1:0] write_burst_packed_addr_92;
  reg [9-1:0] write_burst_packed_stride_93;
  reg [33-1:0] write_burst_packed_length_94;
  reg write_burst_packed_done_95;
  wire [8-1:0] write_burst_packed_ram_addr_96;
  assign write_burst_packed_ram_addr_96 = write_burst_packed_addr_92 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_97;
  assign write_burst_packed_ram_wdata_97 = _maxi_rdata_sb_0 >> 0;
  assign ram_w16_l512_id10_0_1_addr = ((write_burst_packed_fsm_32 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_addr_96 : 'hx;
  assign ram_w16_l512_id10_0_1_wdata = ((write_burst_packed_fsm_32 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_wdata_97 : 'hx;
  assign ram_w16_l512_id10_0_1_wenable = ((write_burst_packed_fsm_32 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  assign ram_w16_l512_id10_0_1_enable = ((write_burst_packed_fsm_32 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  wire [8-1:0] write_burst_packed_ram_addr_98;
  assign write_burst_packed_ram_addr_98 = write_burst_packed_addr_92 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_99;
  assign write_burst_packed_ram_wdata_99 = _maxi_rdata_sb_0 >> 16;
  assign ram_w16_l512_id10_1_1_addr = ((write_burst_packed_fsm_32 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_addr_98 : 'hx;
  assign ram_w16_l512_id10_1_1_wdata = ((write_burst_packed_fsm_32 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_wdata_99 : 'hx;
  assign ram_w16_l512_id10_1_1_wenable = ((write_burst_packed_fsm_32 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  assign ram_w16_l512_id10_1_1_enable = ((write_burst_packed_fsm_32 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  wire [8-1:0] _dma_write_block_high_local_size_100;
  assign _dma_write_block_high_local_size_100 = cparam_conv2d_4_filter_read_size >> 1;
  wire [1-1:0] _dma_write_block_low_local_size_101;
  assign _dma_write_block_low_local_size_101 = cparam_conv2d_4_filter_read_size & { 1{ 1'd1 } };
  wire [8-1:0] _dma_write_block_local_size_102;
  assign _dma_write_block_local_size_102 = (_dma_write_block_low_local_size_101 > 0)? _dma_write_block_high_local_size_100 + 1 : _dma_write_block_high_local_size_100;
  wire [2-1:0] _dma_read_block_high_local_blocksize_103;
  assign _dma_read_block_high_local_blocksize_103 = cparam_conv2d_4_filter_read_block >> 1;
  wire [2-1:0] _dma_read_block_low_local_blocksize_104;
  assign _dma_read_block_low_local_blocksize_104 = cparam_conv2d_4_filter_read_block & { 1{ 1'd1 } };
  wire [2-1:0] _dma_read_block_local_blocksize_105;
  assign _dma_read_block_local_blocksize_105 = (_dma_read_block_low_local_blocksize_104 > 0)? _dma_read_block_high_local_blocksize_103 + 1 : _dma_read_block_high_local_blocksize_103;
  wire [32-1:0] mask_addr_shifted_106;
  assign mask_addr_shifted_106 = conv2d_4_arg_objaddr_1 + conv2d_4_filter_base_offset + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_107;
  assign mask_addr_masked_107 = mask_addr_shifted_106 << 2;
  wire write_burst_block_ram_wvalid_108;
  wire write_burst_block_ram_wquit_109;
  reg [32-1:0] write_burst_packed_fsm_33;
  localparam write_burst_packed_fsm_33_init = 0;
  reg [9-1:0] write_burst_packed_addr_110;
  reg [9-1:0] write_burst_packed_stride_111;
  reg [33-1:0] write_burst_packed_length_112;
  reg write_burst_packed_done_113;
  wire [8-1:0] write_burst_packed_ram_addr_114;
  assign write_burst_packed_ram_addr_114 = write_burst_packed_addr_110 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_115;
  assign write_burst_packed_ram_wdata_115 = _maxi_rdata_sb_0 >> 0;
  assign ram_w16_l512_id0_0_1_wdata = ((write_burst_packed_fsm_33 == 1) && write_burst_block_ram_wvalid_108)? write_burst_packed_ram_wdata_115 : 'hx;
  assign ram_w16_l512_id0_0_1_wenable = ((write_burst_packed_fsm_33 == 1) && write_burst_block_ram_wvalid_108)? 1'd1 : 0;
  wire [8-1:0] write_burst_packed_ram_addr_116;
  assign write_burst_packed_ram_addr_116 = write_burst_packed_addr_110 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_117;
  assign write_burst_packed_ram_wdata_117 = _maxi_rdata_sb_0 >> 16;
  assign ram_w16_l512_id0_1_1_wdata = ((write_burst_packed_fsm_33 == 1) && write_burst_block_ram_wvalid_108)? write_burst_packed_ram_wdata_117 : 'hx;
  assign ram_w16_l512_id0_1_1_wenable = ((write_burst_packed_fsm_33 == 1) && write_burst_block_ram_wvalid_108)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_118;
  wire write_burst_block_ram_wquit_119;
  reg [32-1:0] write_burst_packed_fsm_34;
  localparam write_burst_packed_fsm_34_init = 0;
  reg [9-1:0] write_burst_packed_addr_120;
  reg [9-1:0] write_burst_packed_stride_121;
  reg [33-1:0] write_burst_packed_length_122;
  reg write_burst_packed_done_123;
  wire [8-1:0] write_burst_packed_ram_addr_124;
  assign write_burst_packed_ram_addr_124 = write_burst_packed_addr_120 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_125;
  assign write_burst_packed_ram_wdata_125 = _maxi_rdata_sb_0 >> 0;
  wire [8-1:0] write_burst_packed_ram_addr_126;
  assign write_burst_packed_ram_addr_126 = write_burst_packed_addr_120 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_127;
  assign write_burst_packed_ram_wdata_127 = _maxi_rdata_sb_0 >> 16;
  wire write_burst_block_ram_wvalid_128;
  wire write_burst_block_ram_wquit_129;
  reg [32-1:0] write_burst_packed_fsm_35;
  localparam write_burst_packed_fsm_35_init = 0;
  reg [9-1:0] write_burst_packed_addr_130;
  reg [9-1:0] write_burst_packed_stride_131;
  reg [33-1:0] write_burst_packed_length_132;
  reg write_burst_packed_done_133;
  wire [8-1:0] write_burst_packed_ram_addr_134;
  assign write_burst_packed_ram_addr_134 = write_burst_packed_addr_130 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_135;
  assign write_burst_packed_ram_wdata_135 = _maxi_rdata_sb_0 >> 0;
  wire [8-1:0] write_burst_packed_ram_addr_136;
  assign write_burst_packed_ram_addr_136 = write_burst_packed_addr_130 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_137;
  assign write_burst_packed_ram_wdata_137 = _maxi_rdata_sb_0 >> 16;
  wire write_burst_block_ram_wvalid_138;
  wire write_burst_block_ram_wquit_139;
  reg [32-1:0] write_burst_packed_fsm_36;
  localparam write_burst_packed_fsm_36_init = 0;
  reg [9-1:0] write_burst_packed_addr_140;
  reg [9-1:0] write_burst_packed_stride_141;
  reg [33-1:0] write_burst_packed_length_142;
  reg write_burst_packed_done_143;
  wire [8-1:0] write_burst_packed_ram_addr_144;
  assign write_burst_packed_ram_addr_144 = write_burst_packed_addr_140 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_145;
  assign write_burst_packed_ram_wdata_145 = _maxi_rdata_sb_0 >> 0;
  assign ram_w16_l512_id3_0_1_addr = ((write_burst_packed_fsm_36 == 1) && write_burst_block_ram_wvalid_138)? write_burst_packed_ram_addr_144 : 'hx;
  assign ram_w16_l512_id3_0_1_wdata = ((write_burst_packed_fsm_36 == 1) && write_burst_block_ram_wvalid_138)? write_burst_packed_ram_wdata_145 : 'hx;
  assign ram_w16_l512_id3_0_1_wenable = ((write_burst_packed_fsm_36 == 1) && write_burst_block_ram_wvalid_138)? 1'd1 : 0;
  assign ram_w16_l512_id3_0_1_enable = ((write_burst_packed_fsm_36 == 1) && write_burst_block_ram_wvalid_138)? 1'd1 : 0;
  wire [8-1:0] write_burst_packed_ram_addr_146;
  assign write_burst_packed_ram_addr_146 = write_burst_packed_addr_140 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_147;
  assign write_burst_packed_ram_wdata_147 = _maxi_rdata_sb_0 >> 16;
  assign ram_w16_l512_id3_1_1_addr = ((write_burst_packed_fsm_36 == 1) && write_burst_block_ram_wvalid_138)? write_burst_packed_ram_addr_146 : 'hx;
  assign ram_w16_l512_id3_1_1_wdata = ((write_burst_packed_fsm_36 == 1) && write_burst_block_ram_wvalid_138)? write_burst_packed_ram_wdata_147 : 'hx;
  assign ram_w16_l512_id3_1_1_wenable = ((write_burst_packed_fsm_36 == 1) && write_burst_block_ram_wvalid_138)? 1'd1 : 0;
  assign ram_w16_l512_id3_1_1_enable = ((write_burst_packed_fsm_36 == 1) && write_burst_block_ram_wvalid_138)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_148;
  wire write_burst_block_ram_wquit_149;
  reg [32-1:0] write_burst_packed_fsm_37;
  localparam write_burst_packed_fsm_37_init = 0;
  reg [9-1:0] write_burst_packed_addr_150;
  reg [9-1:0] write_burst_packed_stride_151;
  reg [33-1:0] write_burst_packed_length_152;
  reg write_burst_packed_done_153;
  wire [8-1:0] write_burst_packed_ram_addr_154;
  assign write_burst_packed_ram_addr_154 = write_burst_packed_addr_150 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_155;
  assign write_burst_packed_ram_wdata_155 = _maxi_rdata_sb_0 >> 0;
  assign ram_w16_l512_id4_0_1_addr = ((write_burst_packed_fsm_37 == 1) && write_burst_block_ram_wvalid_148)? write_burst_packed_ram_addr_154 : 'hx;
  assign ram_w16_l512_id4_0_1_wdata = ((write_burst_packed_fsm_37 == 1) && write_burst_block_ram_wvalid_148)? write_burst_packed_ram_wdata_155 : 'hx;
  assign ram_w16_l512_id4_0_1_wenable = ((write_burst_packed_fsm_37 == 1) && write_burst_block_ram_wvalid_148)? 1'd1 : 0;
  assign ram_w16_l512_id4_0_1_enable = ((write_burst_packed_fsm_37 == 1) && write_burst_block_ram_wvalid_148)? 1'd1 : 0;
  wire [8-1:0] write_burst_packed_ram_addr_156;
  assign write_burst_packed_ram_addr_156 = write_burst_packed_addr_150 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_157;
  assign write_burst_packed_ram_wdata_157 = _maxi_rdata_sb_0 >> 16;
  assign ram_w16_l512_id4_1_1_addr = ((write_burst_packed_fsm_37 == 1) && write_burst_block_ram_wvalid_148)? write_burst_packed_ram_addr_156 : 'hx;
  assign ram_w16_l512_id4_1_1_wdata = ((write_burst_packed_fsm_37 == 1) && write_burst_block_ram_wvalid_148)? write_burst_packed_ram_wdata_157 : 'hx;
  assign ram_w16_l512_id4_1_1_wenable = ((write_burst_packed_fsm_37 == 1) && write_burst_block_ram_wvalid_148)? 1'd1 : 0;
  assign ram_w16_l512_id4_1_1_enable = ((write_burst_packed_fsm_37 == 1) && write_burst_block_ram_wvalid_148)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_158;
  wire write_burst_block_ram_wquit_159;
  reg [32-1:0] write_burst_packed_fsm_38;
  localparam write_burst_packed_fsm_38_init = 0;
  reg [9-1:0] write_burst_packed_addr_160;
  reg [9-1:0] write_burst_packed_stride_161;
  reg [33-1:0] write_burst_packed_length_162;
  reg write_burst_packed_done_163;
  wire [8-1:0] write_burst_packed_ram_addr_164;
  assign write_burst_packed_ram_addr_164 = write_burst_packed_addr_160 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_165;
  assign write_burst_packed_ram_wdata_165 = _maxi_rdata_sb_0 >> 0;
  assign ram_w16_l512_id5_0_1_addr = ((write_burst_packed_fsm_38 == 1) && write_burst_block_ram_wvalid_158)? write_burst_packed_ram_addr_164 : 'hx;
  assign ram_w16_l512_id5_0_1_wdata = ((write_burst_packed_fsm_38 == 1) && write_burst_block_ram_wvalid_158)? write_burst_packed_ram_wdata_165 : 'hx;
  assign ram_w16_l512_id5_0_1_wenable = ((write_burst_packed_fsm_38 == 1) && write_burst_block_ram_wvalid_158)? 1'd1 : 0;
  assign ram_w16_l512_id5_0_1_enable = ((write_burst_packed_fsm_38 == 1) && write_burst_block_ram_wvalid_158)? 1'd1 : 0;
  wire [8-1:0] write_burst_packed_ram_addr_166;
  assign write_burst_packed_ram_addr_166 = write_burst_packed_addr_160 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_167;
  assign write_burst_packed_ram_wdata_167 = _maxi_rdata_sb_0 >> 16;
  assign ram_w16_l512_id5_1_1_addr = ((write_burst_packed_fsm_38 == 1) && write_burst_block_ram_wvalid_158)? write_burst_packed_ram_addr_166 : 'hx;
  assign ram_w16_l512_id5_1_1_wdata = ((write_burst_packed_fsm_38 == 1) && write_burst_block_ram_wvalid_158)? write_burst_packed_ram_wdata_167 : 'hx;
  assign ram_w16_l512_id5_1_1_wenable = ((write_burst_packed_fsm_38 == 1) && write_burst_block_ram_wvalid_158)? 1'd1 : 0;
  assign ram_w16_l512_id5_1_1_enable = ((write_burst_packed_fsm_38 == 1) && write_burst_block_ram_wvalid_158)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_168;
  wire write_burst_block_ram_wquit_169;
  reg [32-1:0] write_burst_packed_fsm_39;
  localparam write_burst_packed_fsm_39_init = 0;
  reg [9-1:0] write_burst_packed_addr_170;
  reg [9-1:0] write_burst_packed_stride_171;
  reg [33-1:0] write_burst_packed_length_172;
  reg write_burst_packed_done_173;
  wire [8-1:0] write_burst_packed_ram_addr_174;
  assign write_burst_packed_ram_addr_174 = write_burst_packed_addr_170 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_175;
  assign write_burst_packed_ram_wdata_175 = _maxi_rdata_sb_0 >> 0;
  assign ram_w16_l512_id6_0_1_addr = ((write_burst_packed_fsm_39 == 1) && write_burst_block_ram_wvalid_168)? write_burst_packed_ram_addr_174 : 'hx;
  assign ram_w16_l512_id6_0_1_wdata = ((write_burst_packed_fsm_39 == 1) && write_burst_block_ram_wvalid_168)? write_burst_packed_ram_wdata_175 : 'hx;
  assign ram_w16_l512_id6_0_1_wenable = ((write_burst_packed_fsm_39 == 1) && write_burst_block_ram_wvalid_168)? 1'd1 : 0;
  assign ram_w16_l512_id6_0_1_enable = ((write_burst_packed_fsm_39 == 1) && write_burst_block_ram_wvalid_168)? 1'd1 : 0;
  wire [8-1:0] write_burst_packed_ram_addr_176;
  assign write_burst_packed_ram_addr_176 = write_burst_packed_addr_170 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_177;
  assign write_burst_packed_ram_wdata_177 = _maxi_rdata_sb_0 >> 16;
  assign ram_w16_l512_id6_1_1_addr = ((write_burst_packed_fsm_39 == 1) && write_burst_block_ram_wvalid_168)? write_burst_packed_ram_addr_176 : 'hx;
  assign ram_w16_l512_id6_1_1_wdata = ((write_burst_packed_fsm_39 == 1) && write_burst_block_ram_wvalid_168)? write_burst_packed_ram_wdata_177 : 'hx;
  assign ram_w16_l512_id6_1_1_wenable = ((write_burst_packed_fsm_39 == 1) && write_burst_block_ram_wvalid_168)? 1'd1 : 0;
  assign ram_w16_l512_id6_1_1_enable = ((write_burst_packed_fsm_39 == 1) && write_burst_block_ram_wvalid_168)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_178;
  wire write_burst_block_ram_wquit_179;
  reg [32-1:0] write_burst_packed_fsm_40;
  localparam write_burst_packed_fsm_40_init = 0;
  reg [9-1:0] write_burst_packed_addr_180;
  reg [9-1:0] write_burst_packed_stride_181;
  reg [33-1:0] write_burst_packed_length_182;
  reg write_burst_packed_done_183;
  wire [8-1:0] write_burst_packed_ram_addr_184;
  assign write_burst_packed_ram_addr_184 = write_burst_packed_addr_180 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_185;
  assign write_burst_packed_ram_wdata_185 = _maxi_rdata_sb_0 >> 0;
  assign ram_w16_l512_id7_0_1_addr = ((write_burst_packed_fsm_40 == 1) && write_burst_block_ram_wvalid_178)? write_burst_packed_ram_addr_184 : 'hx;
  assign ram_w16_l512_id7_0_1_wdata = ((write_burst_packed_fsm_40 == 1) && write_burst_block_ram_wvalid_178)? write_burst_packed_ram_wdata_185 : 'hx;
  assign ram_w16_l512_id7_0_1_wenable = ((write_burst_packed_fsm_40 == 1) && write_burst_block_ram_wvalid_178)? 1'd1 : 0;
  assign ram_w16_l512_id7_0_1_enable = ((write_burst_packed_fsm_40 == 1) && write_burst_block_ram_wvalid_178)? 1'd1 : 0;
  wire [8-1:0] write_burst_packed_ram_addr_186;
  assign write_burst_packed_ram_addr_186 = write_burst_packed_addr_180 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_187;
  assign write_burst_packed_ram_wdata_187 = _maxi_rdata_sb_0 >> 16;
  assign ram_w16_l512_id7_1_1_addr = ((write_burst_packed_fsm_40 == 1) && write_burst_block_ram_wvalid_178)? write_burst_packed_ram_addr_186 : 'hx;
  assign ram_w16_l512_id7_1_1_wdata = ((write_burst_packed_fsm_40 == 1) && write_burst_block_ram_wvalid_178)? write_burst_packed_ram_wdata_187 : 'hx;
  assign ram_w16_l512_id7_1_1_wenable = ((write_burst_packed_fsm_40 == 1) && write_burst_block_ram_wvalid_178)? 1'd1 : 0;
  assign ram_w16_l512_id7_1_1_enable = ((write_burst_packed_fsm_40 == 1) && write_burst_block_ram_wvalid_178)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_188;
  wire write_burst_block_ram_wquit_189;
  reg [32-1:0] write_burst_packed_fsm_41;
  localparam write_burst_packed_fsm_41_init = 0;
  reg [9-1:0] write_burst_packed_addr_190;
  reg [9-1:0] write_burst_packed_stride_191;
  reg [33-1:0] write_burst_packed_length_192;
  reg write_burst_packed_done_193;
  wire [8-1:0] write_burst_packed_ram_addr_194;
  assign write_burst_packed_ram_addr_194 = write_burst_packed_addr_190 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_195;
  assign write_burst_packed_ram_wdata_195 = _maxi_rdata_sb_0 >> 0;
  assign ram_w16_l512_id8_0_1_addr = ((write_burst_packed_fsm_41 == 1) && write_burst_block_ram_wvalid_188)? write_burst_packed_ram_addr_194 : 'hx;
  assign ram_w16_l512_id8_0_1_wdata = ((write_burst_packed_fsm_41 == 1) && write_burst_block_ram_wvalid_188)? write_burst_packed_ram_wdata_195 : 'hx;
  assign ram_w16_l512_id8_0_1_wenable = ((write_burst_packed_fsm_41 == 1) && write_burst_block_ram_wvalid_188)? 1'd1 : 0;
  assign ram_w16_l512_id8_0_1_enable = ((write_burst_packed_fsm_41 == 1) && write_burst_block_ram_wvalid_188)? 1'd1 : 0;
  wire [8-1:0] write_burst_packed_ram_addr_196;
  assign write_burst_packed_ram_addr_196 = write_burst_packed_addr_190 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_197;
  assign write_burst_packed_ram_wdata_197 = _maxi_rdata_sb_0 >> 16;
  assign ram_w16_l512_id8_1_1_addr = ((write_burst_packed_fsm_41 == 1) && write_burst_block_ram_wvalid_188)? write_burst_packed_ram_addr_196 : 'hx;
  assign ram_w16_l512_id8_1_1_wdata = ((write_burst_packed_fsm_41 == 1) && write_burst_block_ram_wvalid_188)? write_burst_packed_ram_wdata_197 : 'hx;
  assign ram_w16_l512_id8_1_1_wenable = ((write_burst_packed_fsm_41 == 1) && write_burst_block_ram_wvalid_188)? 1'd1 : 0;
  assign ram_w16_l512_id8_1_1_enable = ((write_burst_packed_fsm_41 == 1) && write_burst_block_ram_wvalid_188)? 1'd1 : 0;
  reg [32-1:0] write_burst_block_fsm_42;
  localparam write_burst_block_fsm_42_init = 0;
  reg [33-1:0] write_burst_block_length_198;
  reg [32-1:0] write_burst_block_blocksize_199;
  reg write_burst_block_done_200;
  reg [32-1:0] write_burst_block_count_201;
  assign write_burst_block_ram_wvalid_108 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_42 == 1);
  assign write_burst_block_ram_wquit_109 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1);
  assign write_burst_block_ram_wvalid_118 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_42 == 2);
  assign write_burst_block_ram_wquit_119 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1);
  assign write_burst_block_ram_wvalid_128 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_42 == 3);
  assign write_burst_block_ram_wquit_129 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1);
  assign write_burst_block_ram_wvalid_138 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_42 == 4);
  assign write_burst_block_ram_wquit_139 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1);
  assign write_burst_block_ram_wvalid_148 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_42 == 5);
  assign write_burst_block_ram_wquit_149 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1);
  assign write_burst_block_ram_wvalid_158 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_42 == 6);
  assign write_burst_block_ram_wquit_159 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1);
  assign write_burst_block_ram_wvalid_168 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_42 == 7);
  assign write_burst_block_ram_wquit_169 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1);
  assign write_burst_block_ram_wvalid_178 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_42 == 8);
  assign write_burst_block_ram_wquit_179 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1);
  assign write_burst_block_ram_wvalid_188 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_42 == 9);
  assign write_burst_block_ram_wquit_189 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1);
  wire [32-1:0] conv2d_4_mux_act_gaddr_0;
  assign conv2d_4_mux_act_gaddr_0 = (conv2d_4_row_select == 0)? conv2d_4_arg_objaddr_0 + (conv2d_4_act_base_offset + cparam_conv2d_4_act_offset_values_0) : 
                                    (conv2d_4_row_select == 1)? conv2d_4_arg_objaddr_0 + (conv2d_4_act_base_offset + cparam_conv2d_4_act_offset_values_2) : 
                                    (conv2d_4_row_select == 2)? conv2d_4_arg_objaddr_0 + (conv2d_4_act_base_offset + cparam_conv2d_4_act_offset_values_1) : 1'd0;
  wire [32-1:0] conv2d_4_mux_act_gaddr_1;
  assign conv2d_4_mux_act_gaddr_1 = (conv2d_4_row_select == 0)? conv2d_4_arg_objaddr_0 + (conv2d_4_act_base_offset + cparam_conv2d_4_act_offset_values_1) : 
                                    (conv2d_4_row_select == 1)? conv2d_4_arg_objaddr_0 + (conv2d_4_act_base_offset + cparam_conv2d_4_act_offset_values_0) : 
                                    (conv2d_4_row_select == 2)? conv2d_4_arg_objaddr_0 + (conv2d_4_act_base_offset + cparam_conv2d_4_act_offset_values_2) : 1'd0;
  wire [32-1:0] conv2d_4_mux_act_gaddr_2;
  assign conv2d_4_mux_act_gaddr_2 = (conv2d_4_row_select == 0)? conv2d_4_arg_objaddr_0 + (conv2d_4_act_base_offset + cparam_conv2d_4_act_offset_values_2) : 
                                    (conv2d_4_row_select == 1)? conv2d_4_arg_objaddr_0 + (conv2d_4_act_base_offset + cparam_conv2d_4_act_offset_values_1) : 
                                    (conv2d_4_row_select == 2)? conv2d_4_arg_objaddr_0 + (conv2d_4_act_base_offset + cparam_conv2d_4_act_offset_values_0) : 1'd0;
  wire conv2d_4_dma_pad_mask_0;
  assign conv2d_4_dma_pad_mask_0 = (conv2d_4_row_count + 0 < cparam_conv2d_4_pad_row_top) || (conv2d_4_row_count + 0 >= cparam_conv2d_4_act_num_row + cparam_conv2d_4_pad_row_top);
  wire conv2d_4_dma_pad_mask_1;
  assign conv2d_4_dma_pad_mask_1 = (conv2d_4_row_count + 1 < cparam_conv2d_4_pad_row_top) || (conv2d_4_row_count + 1 >= cparam_conv2d_4_act_num_row + cparam_conv2d_4_pad_row_top);
  wire conv2d_4_dma_pad_mask_2;
  assign conv2d_4_dma_pad_mask_2 = (conv2d_4_row_count + 2 < cparam_conv2d_4_pad_row_top) || (conv2d_4_row_count + 2 >= cparam_conv2d_4_act_num_row + cparam_conv2d_4_pad_row_top);
  wire conv2d_4_mux_dma_pad_mask_0;
  assign conv2d_4_mux_dma_pad_mask_0 = (conv2d_4_row_select == 0)? conv2d_4_dma_pad_mask_0 : 
                                       (conv2d_4_row_select == 1)? conv2d_4_dma_pad_mask_2 : 
                                       (conv2d_4_row_select == 2)? conv2d_4_dma_pad_mask_1 : 1'd0;
  wire conv2d_4_mux_dma_pad_mask_1;
  assign conv2d_4_mux_dma_pad_mask_1 = (conv2d_4_row_select == 0)? conv2d_4_dma_pad_mask_1 : 
                                       (conv2d_4_row_select == 1)? conv2d_4_dma_pad_mask_0 : 
                                       (conv2d_4_row_select == 2)? conv2d_4_dma_pad_mask_2 : 1'd0;
  wire conv2d_4_mux_dma_pad_mask_2;
  assign conv2d_4_mux_dma_pad_mask_2 = (conv2d_4_row_select == 0)? conv2d_4_dma_pad_mask_2 : 
                                       (conv2d_4_row_select == 1)? conv2d_4_dma_pad_mask_1 : 
                                       (conv2d_4_row_select == 2)? conv2d_4_dma_pad_mask_0 : 1'd0;
  wire conv2d_4_mux_dma_flag_0;
  assign conv2d_4_mux_dma_flag_0 = (conv2d_4_prev_row_select == 0)? conv2d_4_dma_flag_0 : 
                                   (conv2d_4_prev_row_select == 1)? conv2d_4_dma_flag_2 : 
                                   (conv2d_4_prev_row_select == 2)? conv2d_4_dma_flag_1 : 1'd0;
  wire conv2d_4_mux_dma_flag_1;
  assign conv2d_4_mux_dma_flag_1 = (conv2d_4_prev_row_select == 0)? conv2d_4_dma_flag_1 : 
                                   (conv2d_4_prev_row_select == 1)? conv2d_4_dma_flag_0 : 
                                   (conv2d_4_prev_row_select == 2)? conv2d_4_dma_flag_2 : 1'd0;
  wire conv2d_4_mux_dma_flag_2;
  assign conv2d_4_mux_dma_flag_2 = (conv2d_4_prev_row_select == 0)? conv2d_4_dma_flag_2 : 
                                   (conv2d_4_prev_row_select == 1)? conv2d_4_dma_flag_1 : 
                                   (conv2d_4_prev_row_select == 2)? conv2d_4_dma_flag_0 : 1'd0;
  wire [6-1:0] _dma_write_block_high_local_size_202;
  assign _dma_write_block_high_local_size_202 = cparam_conv2d_4_act_read_size >> 1;
  wire [1-1:0] _dma_write_block_low_local_size_203;
  assign _dma_write_block_low_local_size_203 = cparam_conv2d_4_act_read_size & { 1{ 1'd1 } };
  wire [6-1:0] _dma_write_block_local_size_204;
  assign _dma_write_block_local_size_204 = (_dma_write_block_low_local_size_203 > 0)? _dma_write_block_high_local_size_202 + 1 : _dma_write_block_high_local_size_202;
  wire [2-1:0] _dma_read_block_high_local_blocksize_205;
  assign _dma_read_block_high_local_blocksize_205 = cparam_conv2d_4_act_read_block >> 1;
  wire [2-1:0] _dma_read_block_low_local_blocksize_206;
  assign _dma_read_block_low_local_blocksize_206 = cparam_conv2d_4_act_read_block & { 1{ 1'd1 } };
  wire [2-1:0] _dma_read_block_local_blocksize_207;
  assign _dma_read_block_local_blocksize_207 = (_dma_read_block_low_local_blocksize_206 > 0)? _dma_read_block_high_local_blocksize_205 + 1 : _dma_read_block_high_local_blocksize_205;
  wire [32-1:0] mask_addr_shifted_208;
  assign mask_addr_shifted_208 = conv2d_4_mux_act_gaddr_0 + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_209;
  assign mask_addr_masked_209 = mask_addr_shifted_208 << 2;
  wire write_burst_block_ram_wvalid_210;
  wire write_burst_block_ram_wquit_211;
  reg [32-1:0] write_burst_packed_fsm_43;
  localparam write_burst_packed_fsm_43_init = 0;
  reg [9-1:0] write_burst_packed_addr_212;
  reg [9-1:0] write_burst_packed_stride_213;
  reg [33-1:0] write_burst_packed_length_214;
  reg write_burst_packed_done_215;
  wire [8-1:0] write_burst_packed_ram_addr_216;
  assign write_burst_packed_ram_addr_216 = write_burst_packed_addr_212 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_217;
  assign write_burst_packed_ram_wdata_217 = _maxi_rdata_sb_0 >> 0;
  assign ram_w16_l512_id11_0_1_addr = ((write_burst_packed_fsm_43 == 1) && write_burst_block_ram_wvalid_210)? write_burst_packed_ram_addr_216 : 'hx;
  assign ram_w16_l512_id11_0_1_wdata = ((write_burst_packed_fsm_43 == 1) && write_burst_block_ram_wvalid_210)? write_burst_packed_ram_wdata_217 : 'hx;
  assign ram_w16_l512_id11_0_1_wenable = ((write_burst_packed_fsm_43 == 1) && write_burst_block_ram_wvalid_210)? 1'd1 : 0;
  assign ram_w16_l512_id11_0_1_enable = ((write_burst_packed_fsm_43 == 1) && write_burst_block_ram_wvalid_210)? 1'd1 : 0;
  wire [8-1:0] write_burst_packed_ram_addr_218;
  assign write_burst_packed_ram_addr_218 = write_burst_packed_addr_212 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_219;
  assign write_burst_packed_ram_wdata_219 = _maxi_rdata_sb_0 >> 16;
  assign ram_w16_l512_id11_1_1_addr = ((write_burst_packed_fsm_43 == 1) && write_burst_block_ram_wvalid_210)? write_burst_packed_ram_addr_218 : 'hx;
  assign ram_w16_l512_id11_1_1_wdata = ((write_burst_packed_fsm_43 == 1) && write_burst_block_ram_wvalid_210)? write_burst_packed_ram_wdata_219 : 'hx;
  assign ram_w16_l512_id11_1_1_wenable = ((write_burst_packed_fsm_43 == 1) && write_burst_block_ram_wvalid_210)? 1'd1 : 0;
  assign ram_w16_l512_id11_1_1_enable = ((write_burst_packed_fsm_43 == 1) && write_burst_block_ram_wvalid_210)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_220;
  wire write_burst_block_ram_wquit_221;
  reg [32-1:0] write_burst_packed_fsm_44;
  localparam write_burst_packed_fsm_44_init = 0;
  reg [9-1:0] write_burst_packed_addr_222;
  reg [9-1:0] write_burst_packed_stride_223;
  reg [33-1:0] write_burst_packed_length_224;
  reg write_burst_packed_done_225;
  wire [8-1:0] write_burst_packed_ram_addr_226;
  assign write_burst_packed_ram_addr_226 = write_burst_packed_addr_222 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_227;
  assign write_burst_packed_ram_wdata_227 = _maxi_rdata_sb_0 >> 0;
  assign ram_w16_l512_id12_0_1_addr = ((write_burst_packed_fsm_44 == 1) && write_burst_block_ram_wvalid_220)? write_burst_packed_ram_addr_226 : 'hx;
  assign ram_w16_l512_id12_0_1_wdata = ((write_burst_packed_fsm_44 == 1) && write_burst_block_ram_wvalid_220)? write_burst_packed_ram_wdata_227 : 'hx;
  assign ram_w16_l512_id12_0_1_wenable = ((write_burst_packed_fsm_44 == 1) && write_burst_block_ram_wvalid_220)? 1'd1 : 0;
  assign ram_w16_l512_id12_0_1_enable = ((write_burst_packed_fsm_44 == 1) && write_burst_block_ram_wvalid_220)? 1'd1 : 0;
  wire [8-1:0] write_burst_packed_ram_addr_228;
  assign write_burst_packed_ram_addr_228 = write_burst_packed_addr_222 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_229;
  assign write_burst_packed_ram_wdata_229 = _maxi_rdata_sb_0 >> 16;
  assign ram_w16_l512_id12_1_1_addr = ((write_burst_packed_fsm_44 == 1) && write_burst_block_ram_wvalid_220)? write_burst_packed_ram_addr_228 : 'hx;
  assign ram_w16_l512_id12_1_1_wdata = ((write_burst_packed_fsm_44 == 1) && write_burst_block_ram_wvalid_220)? write_burst_packed_ram_wdata_229 : 'hx;
  assign ram_w16_l512_id12_1_1_wenable = ((write_burst_packed_fsm_44 == 1) && write_burst_block_ram_wvalid_220)? 1'd1 : 0;
  assign ram_w16_l512_id12_1_1_enable = ((write_burst_packed_fsm_44 == 1) && write_burst_block_ram_wvalid_220)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_230;
  wire write_burst_block_ram_wquit_231;
  reg [32-1:0] write_burst_packed_fsm_45;
  localparam write_burst_packed_fsm_45_init = 0;
  reg [9-1:0] write_burst_packed_addr_232;
  reg [9-1:0] write_burst_packed_stride_233;
  reg [33-1:0] write_burst_packed_length_234;
  reg write_burst_packed_done_235;
  wire [8-1:0] write_burst_packed_ram_addr_236;
  assign write_burst_packed_ram_addr_236 = write_burst_packed_addr_232 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_237;
  assign write_burst_packed_ram_wdata_237 = _maxi_rdata_sb_0 >> 0;
  assign ram_w16_l512_id13_0_1_addr = ((write_burst_packed_fsm_45 == 1) && write_burst_block_ram_wvalid_230)? write_burst_packed_ram_addr_236 : 'hx;
  assign ram_w16_l512_id13_0_1_wdata = ((write_burst_packed_fsm_45 == 1) && write_burst_block_ram_wvalid_230)? write_burst_packed_ram_wdata_237 : 'hx;
  assign ram_w16_l512_id13_0_1_wenable = ((write_burst_packed_fsm_45 == 1) && write_burst_block_ram_wvalid_230)? 1'd1 : 0;
  assign ram_w16_l512_id13_0_1_enable = ((write_burst_packed_fsm_45 == 1) && write_burst_block_ram_wvalid_230)? 1'd1 : 0;
  wire [8-1:0] write_burst_packed_ram_addr_238;
  assign write_burst_packed_ram_addr_238 = write_burst_packed_addr_232 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_239;
  assign write_burst_packed_ram_wdata_239 = _maxi_rdata_sb_0 >> 16;
  assign ram_w16_l512_id13_1_1_addr = ((write_burst_packed_fsm_45 == 1) && write_burst_block_ram_wvalid_230)? write_burst_packed_ram_addr_238 : 'hx;
  assign ram_w16_l512_id13_1_1_wdata = ((write_burst_packed_fsm_45 == 1) && write_burst_block_ram_wvalid_230)? write_burst_packed_ram_wdata_239 : 'hx;
  assign ram_w16_l512_id13_1_1_wenable = ((write_burst_packed_fsm_45 == 1) && write_burst_block_ram_wvalid_230)? 1'd1 : 0;
  assign ram_w16_l512_id13_1_1_enable = ((write_burst_packed_fsm_45 == 1) && write_burst_block_ram_wvalid_230)? 1'd1 : 0;
  reg [32-1:0] write_burst_block_fsm_46;
  localparam write_burst_block_fsm_46_init = 0;
  reg [33-1:0] write_burst_block_length_240;
  reg [32-1:0] write_burst_block_blocksize_241;
  reg write_burst_block_done_242;
  reg [32-1:0] write_burst_block_count_243;
  assign write_burst_block_ram_wvalid_210 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_46 == 1);
  assign write_burst_block_ram_wquit_211 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_240 <= 1);
  assign write_burst_block_ram_wvalid_220 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_46 == 2);
  assign write_burst_block_ram_wquit_221 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_240 <= 1);
  assign write_burst_block_ram_wvalid_230 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_46 == 3);
  assign write_burst_block_ram_wquit_231 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_240 <= 1);
  wire [6-1:0] _dma_write_block_high_local_size_244;
  assign _dma_write_block_high_local_size_244 = cparam_conv2d_4_act_read_size >> 1;
  wire [1-1:0] _dma_write_block_low_local_size_245;
  assign _dma_write_block_low_local_size_245 = cparam_conv2d_4_act_read_size & { 1{ 1'd1 } };
  wire [6-1:0] _dma_write_block_local_size_246;
  assign _dma_write_block_local_size_246 = (_dma_write_block_low_local_size_245 > 0)? _dma_write_block_high_local_size_244 + 1 : _dma_write_block_high_local_size_244;
  wire [2-1:0] _dma_read_block_high_local_blocksize_247;
  assign _dma_read_block_high_local_blocksize_247 = cparam_conv2d_4_act_read_block >> 1;
  wire [2-1:0] _dma_read_block_low_local_blocksize_248;
  assign _dma_read_block_low_local_blocksize_248 = cparam_conv2d_4_act_read_block & { 1{ 1'd1 } };
  wire [2-1:0] _dma_read_block_local_blocksize_249;
  assign _dma_read_block_local_blocksize_249 = (_dma_read_block_low_local_blocksize_248 > 0)? _dma_read_block_high_local_blocksize_247 + 1 : _dma_read_block_high_local_blocksize_247;
  wire [32-1:0] mask_addr_shifted_250;
  assign mask_addr_shifted_250 = conv2d_4_mux_act_gaddr_1 + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_251;
  assign mask_addr_masked_251 = mask_addr_shifted_250 << 2;
  wire write_burst_block_ram_wvalid_252;
  wire write_burst_block_ram_wquit_253;
  reg [32-1:0] write_burst_packed_fsm_47;
  localparam write_burst_packed_fsm_47_init = 0;
  reg [9-1:0] write_burst_packed_addr_254;
  reg [9-1:0] write_burst_packed_stride_255;
  reg [33-1:0] write_burst_packed_length_256;
  reg write_burst_packed_done_257;
  wire [8-1:0] write_burst_packed_ram_addr_258;
  assign write_burst_packed_ram_addr_258 = write_burst_packed_addr_254 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_259;
  assign write_burst_packed_ram_wdata_259 = _maxi_rdata_sb_0 >> 0;
  assign ram_w16_l512_id14_0_1_addr = ((write_burst_packed_fsm_47 == 1) && write_burst_block_ram_wvalid_252)? write_burst_packed_ram_addr_258 : 'hx;
  assign ram_w16_l512_id14_0_1_wdata = ((write_burst_packed_fsm_47 == 1) && write_burst_block_ram_wvalid_252)? write_burst_packed_ram_wdata_259 : 'hx;
  assign ram_w16_l512_id14_0_1_wenable = ((write_burst_packed_fsm_47 == 1) && write_burst_block_ram_wvalid_252)? 1'd1 : 0;
  assign ram_w16_l512_id14_0_1_enable = ((write_burst_packed_fsm_47 == 1) && write_burst_block_ram_wvalid_252)? 1'd1 : 0;
  wire [8-1:0] write_burst_packed_ram_addr_260;
  assign write_burst_packed_ram_addr_260 = write_burst_packed_addr_254 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_261;
  assign write_burst_packed_ram_wdata_261 = _maxi_rdata_sb_0 >> 16;
  assign ram_w16_l512_id14_1_1_addr = ((write_burst_packed_fsm_47 == 1) && write_burst_block_ram_wvalid_252)? write_burst_packed_ram_addr_260 : 'hx;
  assign ram_w16_l512_id14_1_1_wdata = ((write_burst_packed_fsm_47 == 1) && write_burst_block_ram_wvalid_252)? write_burst_packed_ram_wdata_261 : 'hx;
  assign ram_w16_l512_id14_1_1_wenable = ((write_burst_packed_fsm_47 == 1) && write_burst_block_ram_wvalid_252)? 1'd1 : 0;
  assign ram_w16_l512_id14_1_1_enable = ((write_burst_packed_fsm_47 == 1) && write_burst_block_ram_wvalid_252)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_262;
  wire write_burst_block_ram_wquit_263;
  reg [32-1:0] write_burst_packed_fsm_48;
  localparam write_burst_packed_fsm_48_init = 0;
  reg [9-1:0] write_burst_packed_addr_264;
  reg [9-1:0] write_burst_packed_stride_265;
  reg [33-1:0] write_burst_packed_length_266;
  reg write_burst_packed_done_267;
  wire [8-1:0] write_burst_packed_ram_addr_268;
  assign write_burst_packed_ram_addr_268 = write_burst_packed_addr_264 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_269;
  assign write_burst_packed_ram_wdata_269 = _maxi_rdata_sb_0 >> 0;
  assign ram_w16_l512_id15_0_1_addr = ((write_burst_packed_fsm_48 == 1) && write_burst_block_ram_wvalid_262)? write_burst_packed_ram_addr_268 : 'hx;
  assign ram_w16_l512_id15_0_1_wdata = ((write_burst_packed_fsm_48 == 1) && write_burst_block_ram_wvalid_262)? write_burst_packed_ram_wdata_269 : 'hx;
  assign ram_w16_l512_id15_0_1_wenable = ((write_burst_packed_fsm_48 == 1) && write_burst_block_ram_wvalid_262)? 1'd1 : 0;
  assign ram_w16_l512_id15_0_1_enable = ((write_burst_packed_fsm_48 == 1) && write_burst_block_ram_wvalid_262)? 1'd1 : 0;
  wire [8-1:0] write_burst_packed_ram_addr_270;
  assign write_burst_packed_ram_addr_270 = write_burst_packed_addr_264 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_271;
  assign write_burst_packed_ram_wdata_271 = _maxi_rdata_sb_0 >> 16;
  assign ram_w16_l512_id15_1_1_addr = ((write_burst_packed_fsm_48 == 1) && write_burst_block_ram_wvalid_262)? write_burst_packed_ram_addr_270 : 'hx;
  assign ram_w16_l512_id15_1_1_wdata = ((write_burst_packed_fsm_48 == 1) && write_burst_block_ram_wvalid_262)? write_burst_packed_ram_wdata_271 : 'hx;
  assign ram_w16_l512_id15_1_1_wenable = ((write_burst_packed_fsm_48 == 1) && write_burst_block_ram_wvalid_262)? 1'd1 : 0;
  assign ram_w16_l512_id15_1_1_enable = ((write_burst_packed_fsm_48 == 1) && write_burst_block_ram_wvalid_262)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_272;
  wire write_burst_block_ram_wquit_273;
  reg [32-1:0] write_burst_packed_fsm_49;
  localparam write_burst_packed_fsm_49_init = 0;
  reg [9-1:0] write_burst_packed_addr_274;
  reg [9-1:0] write_burst_packed_stride_275;
  reg [33-1:0] write_burst_packed_length_276;
  reg write_burst_packed_done_277;
  wire [8-1:0] write_burst_packed_ram_addr_278;
  assign write_burst_packed_ram_addr_278 = write_burst_packed_addr_274 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_279;
  assign write_burst_packed_ram_wdata_279 = _maxi_rdata_sb_0 >> 0;
  assign ram_w16_l512_id16_0_1_addr = ((write_burst_packed_fsm_49 == 1) && write_burst_block_ram_wvalid_272)? write_burst_packed_ram_addr_278 : 'hx;
  assign ram_w16_l512_id16_0_1_wdata = ((write_burst_packed_fsm_49 == 1) && write_burst_block_ram_wvalid_272)? write_burst_packed_ram_wdata_279 : 'hx;
  assign ram_w16_l512_id16_0_1_wenable = ((write_burst_packed_fsm_49 == 1) && write_burst_block_ram_wvalid_272)? 1'd1 : 0;
  assign ram_w16_l512_id16_0_1_enable = ((write_burst_packed_fsm_49 == 1) && write_burst_block_ram_wvalid_272)? 1'd1 : 0;
  wire [8-1:0] write_burst_packed_ram_addr_280;
  assign write_burst_packed_ram_addr_280 = write_burst_packed_addr_274 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_281;
  assign write_burst_packed_ram_wdata_281 = _maxi_rdata_sb_0 >> 16;
  assign ram_w16_l512_id16_1_1_addr = ((write_burst_packed_fsm_49 == 1) && write_burst_block_ram_wvalid_272)? write_burst_packed_ram_addr_280 : 'hx;
  assign ram_w16_l512_id16_1_1_wdata = ((write_burst_packed_fsm_49 == 1) && write_burst_block_ram_wvalid_272)? write_burst_packed_ram_wdata_281 : 'hx;
  assign ram_w16_l512_id16_1_1_wenable = ((write_burst_packed_fsm_49 == 1) && write_burst_block_ram_wvalid_272)? 1'd1 : 0;
  assign ram_w16_l512_id16_1_1_enable = ((write_burst_packed_fsm_49 == 1) && write_burst_block_ram_wvalid_272)? 1'd1 : 0;
  reg [32-1:0] write_burst_block_fsm_50;
  localparam write_burst_block_fsm_50_init = 0;
  reg [33-1:0] write_burst_block_length_282;
  reg [32-1:0] write_burst_block_blocksize_283;
  reg write_burst_block_done_284;
  reg [32-1:0] write_burst_block_count_285;
  assign write_burst_block_ram_wvalid_252 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_50 == 1);
  assign write_burst_block_ram_wquit_253 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_282 <= 1);
  assign write_burst_block_ram_wvalid_262 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_50 == 2);
  assign write_burst_block_ram_wquit_263 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_282 <= 1);
  assign write_burst_block_ram_wvalid_272 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_50 == 3);
  assign write_burst_block_ram_wquit_273 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_282 <= 1);
  wire [6-1:0] _dma_write_block_high_local_size_286;
  assign _dma_write_block_high_local_size_286 = cparam_conv2d_4_act_read_size >> 1;
  wire [1-1:0] _dma_write_block_low_local_size_287;
  assign _dma_write_block_low_local_size_287 = cparam_conv2d_4_act_read_size & { 1{ 1'd1 } };
  wire [6-1:0] _dma_write_block_local_size_288;
  assign _dma_write_block_local_size_288 = (_dma_write_block_low_local_size_287 > 0)? _dma_write_block_high_local_size_286 + 1 : _dma_write_block_high_local_size_286;
  wire [2-1:0] _dma_read_block_high_local_blocksize_289;
  assign _dma_read_block_high_local_blocksize_289 = cparam_conv2d_4_act_read_block >> 1;
  wire [2-1:0] _dma_read_block_low_local_blocksize_290;
  assign _dma_read_block_low_local_blocksize_290 = cparam_conv2d_4_act_read_block & { 1{ 1'd1 } };
  wire [2-1:0] _dma_read_block_local_blocksize_291;
  assign _dma_read_block_local_blocksize_291 = (_dma_read_block_low_local_blocksize_290 > 0)? _dma_read_block_high_local_blocksize_289 + 1 : _dma_read_block_high_local_blocksize_289;
  wire [32-1:0] mask_addr_shifted_292;
  assign mask_addr_shifted_292 = conv2d_4_mux_act_gaddr_2 + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_293;
  assign mask_addr_masked_293 = mask_addr_shifted_292 << 2;
  wire write_burst_block_ram_wvalid_294;
  wire write_burst_block_ram_wquit_295;
  reg [32-1:0] write_burst_packed_fsm_51;
  localparam write_burst_packed_fsm_51_init = 0;
  reg [9-1:0] write_burst_packed_addr_296;
  reg [9-1:0] write_burst_packed_stride_297;
  reg [33-1:0] write_burst_packed_length_298;
  reg write_burst_packed_done_299;
  wire [8-1:0] write_burst_packed_ram_addr_300;
  assign write_burst_packed_ram_addr_300 = write_burst_packed_addr_296 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_301;
  assign write_burst_packed_ram_wdata_301 = _maxi_rdata_sb_0 >> 0;
  assign ram_w16_l512_id17_0_1_addr = ((write_burst_packed_fsm_51 == 1) && write_burst_block_ram_wvalid_294)? write_burst_packed_ram_addr_300 : 'hx;
  assign ram_w16_l512_id17_0_1_wdata = ((write_burst_packed_fsm_51 == 1) && write_burst_block_ram_wvalid_294)? write_burst_packed_ram_wdata_301 : 'hx;
  assign ram_w16_l512_id17_0_1_wenable = ((write_burst_packed_fsm_51 == 1) && write_burst_block_ram_wvalid_294)? 1'd1 : 0;
  assign ram_w16_l512_id17_0_1_enable = ((write_burst_packed_fsm_51 == 1) && write_burst_block_ram_wvalid_294)? 1'd1 : 0;
  wire [8-1:0] write_burst_packed_ram_addr_302;
  assign write_burst_packed_ram_addr_302 = write_burst_packed_addr_296 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_303;
  assign write_burst_packed_ram_wdata_303 = _maxi_rdata_sb_0 >> 16;
  assign ram_w16_l512_id17_1_1_addr = ((write_burst_packed_fsm_51 == 1) && write_burst_block_ram_wvalid_294)? write_burst_packed_ram_addr_302 : 'hx;
  assign ram_w16_l512_id17_1_1_wdata = ((write_burst_packed_fsm_51 == 1) && write_burst_block_ram_wvalid_294)? write_burst_packed_ram_wdata_303 : 'hx;
  assign ram_w16_l512_id17_1_1_wenable = ((write_burst_packed_fsm_51 == 1) && write_burst_block_ram_wvalid_294)? 1'd1 : 0;
  assign ram_w16_l512_id17_1_1_enable = ((write_burst_packed_fsm_51 == 1) && write_burst_block_ram_wvalid_294)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_304;
  wire write_burst_block_ram_wquit_305;
  reg [32-1:0] write_burst_packed_fsm_52;
  localparam write_burst_packed_fsm_52_init = 0;
  reg [9-1:0] write_burst_packed_addr_306;
  reg [9-1:0] write_burst_packed_stride_307;
  reg [33-1:0] write_burst_packed_length_308;
  reg write_burst_packed_done_309;
  wire [8-1:0] write_burst_packed_ram_addr_310;
  assign write_burst_packed_ram_addr_310 = write_burst_packed_addr_306 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_311;
  assign write_burst_packed_ram_wdata_311 = _maxi_rdata_sb_0 >> 0;
  assign ram_w16_l512_id18_0_1_addr = ((write_burst_packed_fsm_52 == 1) && write_burst_block_ram_wvalid_304)? write_burst_packed_ram_addr_310 : 'hx;
  assign ram_w16_l512_id18_0_1_wdata = ((write_burst_packed_fsm_52 == 1) && write_burst_block_ram_wvalid_304)? write_burst_packed_ram_wdata_311 : 'hx;
  assign ram_w16_l512_id18_0_1_wenable = ((write_burst_packed_fsm_52 == 1) && write_burst_block_ram_wvalid_304)? 1'd1 : 0;
  assign ram_w16_l512_id18_0_1_enable = ((write_burst_packed_fsm_52 == 1) && write_burst_block_ram_wvalid_304)? 1'd1 : 0;
  wire [8-1:0] write_burst_packed_ram_addr_312;
  assign write_burst_packed_ram_addr_312 = write_burst_packed_addr_306 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_313;
  assign write_burst_packed_ram_wdata_313 = _maxi_rdata_sb_0 >> 16;
  assign ram_w16_l512_id18_1_1_addr = ((write_burst_packed_fsm_52 == 1) && write_burst_block_ram_wvalid_304)? write_burst_packed_ram_addr_312 : 'hx;
  assign ram_w16_l512_id18_1_1_wdata = ((write_burst_packed_fsm_52 == 1) && write_burst_block_ram_wvalid_304)? write_burst_packed_ram_wdata_313 : 'hx;
  assign ram_w16_l512_id18_1_1_wenable = ((write_burst_packed_fsm_52 == 1) && write_burst_block_ram_wvalid_304)? 1'd1 : 0;
  assign ram_w16_l512_id18_1_1_enable = ((write_burst_packed_fsm_52 == 1) && write_burst_block_ram_wvalid_304)? 1'd1 : 0;
  wire write_burst_block_ram_wvalid_314;
  wire write_burst_block_ram_wquit_315;
  reg [32-1:0] write_burst_packed_fsm_53;
  localparam write_burst_packed_fsm_53_init = 0;
  reg [9-1:0] write_burst_packed_addr_316;
  reg [9-1:0] write_burst_packed_stride_317;
  reg [33-1:0] write_burst_packed_length_318;
  reg write_burst_packed_done_319;
  wire [8-1:0] write_burst_packed_ram_addr_320;
  assign write_burst_packed_ram_addr_320 = write_burst_packed_addr_316 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_321;
  assign write_burst_packed_ram_wdata_321 = _maxi_rdata_sb_0 >> 0;
  assign ram_w16_l512_id19_0_1_addr = ((write_burst_packed_fsm_53 == 1) && write_burst_block_ram_wvalid_314)? write_burst_packed_ram_addr_320 : 'hx;
  assign ram_w16_l512_id19_0_1_wdata = ((write_burst_packed_fsm_53 == 1) && write_burst_block_ram_wvalid_314)? write_burst_packed_ram_wdata_321 : 'hx;
  assign ram_w16_l512_id19_0_1_wenable = ((write_burst_packed_fsm_53 == 1) && write_burst_block_ram_wvalid_314)? 1'd1 : 0;
  assign ram_w16_l512_id19_0_1_enable = ((write_burst_packed_fsm_53 == 1) && write_burst_block_ram_wvalid_314)? 1'd1 : 0;
  wire [8-1:0] write_burst_packed_ram_addr_322;
  assign write_burst_packed_ram_addr_322 = write_burst_packed_addr_316 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_323;
  assign write_burst_packed_ram_wdata_323 = _maxi_rdata_sb_0 >> 16;
  assign ram_w16_l512_id19_1_1_addr = ((write_burst_packed_fsm_53 == 1) && write_burst_block_ram_wvalid_314)? write_burst_packed_ram_addr_322 : 'hx;
  assign ram_w16_l512_id19_1_1_wdata = ((write_burst_packed_fsm_53 == 1) && write_burst_block_ram_wvalid_314)? write_burst_packed_ram_wdata_323 : 'hx;
  assign ram_w16_l512_id19_1_1_wenable = ((write_burst_packed_fsm_53 == 1) && write_burst_block_ram_wvalid_314)? 1'd1 : 0;
  assign ram_w16_l512_id19_1_1_enable = ((write_burst_packed_fsm_53 == 1) && write_burst_block_ram_wvalid_314)? 1'd1 : 0;
  reg [32-1:0] write_burst_block_fsm_54;
  localparam write_burst_block_fsm_54_init = 0;
  reg [33-1:0] write_burst_block_length_324;
  reg [32-1:0] write_burst_block_blocksize_325;
  reg write_burst_block_done_326;
  reg [32-1:0] write_burst_block_count_327;
  assign write_burst_block_ram_wvalid_294 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_54 == 1);
  assign write_burst_block_ram_wquit_295 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_324 <= 1);
  assign write_burst_block_ram_wvalid_304 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_54 == 2);
  assign write_burst_block_ram_wquit_305 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_324 <= 1);
  assign write_burst_block_ram_wvalid_314 = _maxi_rvalid_sb_0 && (write_burst_block_fsm_54 == 3);
  assign write_burst_block_ram_wquit_315 = 0 || _maxi_rvalid_sb_0 && 0 || _maxi_rvalid_sb_0 && (write_burst_block_length_324 <= 1);
  reg [32-1:0] conv2d_4_comp_fsm;
  localparam conv2d_4_comp_fsm_init = 0;
  reg [32-1:0] conv2d_4_filter_page_comp_offset_buf;
  reg [32-1:0] conv2d_4_act_page_comp_offset_buf_0;
  reg [32-1:0] conv2d_4_act_page_comp_offset_buf_1;
  reg [32-1:0] conv2d_4_act_page_comp_offset_buf_2;
  reg [32-1:0] conv2d_4_out_page_comp_offset_buf;
  reg [32-1:0] conv2d_4_row_count_buf;
  reg [2-1:0] conv2d_4_row_select_buf;
  reg [32-1:0] conv2d_4_och_count_buf;
  wire conv2d_4_stream_pad_mask_0_0;
  assign conv2d_4_stream_pad_mask_0_0 = (conv2d_4_col_count + 0 < cparam_conv2d_4_pad_col_left) || (conv2d_4_col_count + 0 >= cparam_conv2d_4_act_num_col + cparam_conv2d_4_pad_col_left) || (conv2d_4_row_count_buf + 0 < cparam_conv2d_4_pad_row_top) || (conv2d_4_row_count_buf + 0 >= cparam_conv2d_4_act_num_row + cparam_conv2d_4_pad_row_top);
  wire conv2d_4_stream_pad_mask_0_1;
  assign conv2d_4_stream_pad_mask_0_1 = (conv2d_4_col_count + 1 < cparam_conv2d_4_pad_col_left) || (conv2d_4_col_count + 1 >= cparam_conv2d_4_act_num_col + cparam_conv2d_4_pad_col_left) || (conv2d_4_row_count_buf + 0 < cparam_conv2d_4_pad_row_top) || (conv2d_4_row_count_buf + 0 >= cparam_conv2d_4_act_num_row + cparam_conv2d_4_pad_row_top);
  wire conv2d_4_stream_pad_mask_0_2;
  assign conv2d_4_stream_pad_mask_0_2 = (conv2d_4_col_count + 2 < cparam_conv2d_4_pad_col_left) || (conv2d_4_col_count + 2 >= cparam_conv2d_4_act_num_col + cparam_conv2d_4_pad_col_left) || (conv2d_4_row_count_buf + 0 < cparam_conv2d_4_pad_row_top) || (conv2d_4_row_count_buf + 0 >= cparam_conv2d_4_act_num_row + cparam_conv2d_4_pad_row_top);
  wire conv2d_4_stream_pad_mask_1_0;
  assign conv2d_4_stream_pad_mask_1_0 = (conv2d_4_col_count + 0 < cparam_conv2d_4_pad_col_left) || (conv2d_4_col_count + 0 >= cparam_conv2d_4_act_num_col + cparam_conv2d_4_pad_col_left) || (conv2d_4_row_count_buf + 1 < cparam_conv2d_4_pad_row_top) || (conv2d_4_row_count_buf + 1 >= cparam_conv2d_4_act_num_row + cparam_conv2d_4_pad_row_top);
  wire conv2d_4_stream_pad_mask_1_1;
  assign conv2d_4_stream_pad_mask_1_1 = (conv2d_4_col_count + 1 < cparam_conv2d_4_pad_col_left) || (conv2d_4_col_count + 1 >= cparam_conv2d_4_act_num_col + cparam_conv2d_4_pad_col_left) || (conv2d_4_row_count_buf + 1 < cparam_conv2d_4_pad_row_top) || (conv2d_4_row_count_buf + 1 >= cparam_conv2d_4_act_num_row + cparam_conv2d_4_pad_row_top);
  wire conv2d_4_stream_pad_mask_1_2;
  assign conv2d_4_stream_pad_mask_1_2 = (conv2d_4_col_count + 2 < cparam_conv2d_4_pad_col_left) || (conv2d_4_col_count + 2 >= cparam_conv2d_4_act_num_col + cparam_conv2d_4_pad_col_left) || (conv2d_4_row_count_buf + 1 < cparam_conv2d_4_pad_row_top) || (conv2d_4_row_count_buf + 1 >= cparam_conv2d_4_act_num_row + cparam_conv2d_4_pad_row_top);
  wire conv2d_4_stream_pad_mask_2_0;
  assign conv2d_4_stream_pad_mask_2_0 = (conv2d_4_col_count + 0 < cparam_conv2d_4_pad_col_left) || (conv2d_4_col_count + 0 >= cparam_conv2d_4_act_num_col + cparam_conv2d_4_pad_col_left) || (conv2d_4_row_count_buf + 2 < cparam_conv2d_4_pad_row_top) || (conv2d_4_row_count_buf + 2 >= cparam_conv2d_4_act_num_row + cparam_conv2d_4_pad_row_top);
  wire conv2d_4_stream_pad_mask_2_1;
  assign conv2d_4_stream_pad_mask_2_1 = (conv2d_4_col_count + 1 < cparam_conv2d_4_pad_col_left) || (conv2d_4_col_count + 1 >= cparam_conv2d_4_act_num_col + cparam_conv2d_4_pad_col_left) || (conv2d_4_row_count_buf + 2 < cparam_conv2d_4_pad_row_top) || (conv2d_4_row_count_buf + 2 >= cparam_conv2d_4_act_num_row + cparam_conv2d_4_pad_row_top);
  wire conv2d_4_stream_pad_mask_2_2;
  assign conv2d_4_stream_pad_mask_2_2 = (conv2d_4_col_count + 2 < cparam_conv2d_4_pad_col_left) || (conv2d_4_col_count + 2 >= cparam_conv2d_4_act_num_col + cparam_conv2d_4_pad_col_left) || (conv2d_4_row_count_buf + 2 < cparam_conv2d_4_pad_row_top) || (conv2d_4_row_count_buf + 2 >= cparam_conv2d_4_act_num_row + cparam_conv2d_4_pad_row_top);
  reg [9-1:0] conv2d_4_stream_pad_masks;
  wire [1-1:0] stream_conv2d_4_parameter_0_data;
  wire [2-1:0] stream_conv2d_4_parameter_1_data;
  wire [2-1:0] stream_conv2d_4_parameter_2_data;
  wire [9-1:0] stream_conv2d_4_parameter_3_data;
  wire [1-1:0] stream_conv2d_4_parameter_4_data;
  wire [1-1:0] stream_conv2d_4__reduce_reset_data;
  wire [1-1:0] stream_conv2d_4_parameter_6_data;
  wire [16-1:0] stream_conv2d_4_source_7_data;
  wire [1-1:0] stream_conv2d_4_parameter_8_data;
  wire [16-1:0] stream_conv2d_4_source_9_data;
  wire [1-1:0] stream_conv2d_4_parameter_10_data;
  wire [16-1:0] stream_conv2d_4_source_11_data;
  wire [1-1:0] stream_conv2d_4_parameter_12_data;
  wire [16-1:0] stream_conv2d_4_source_13_data;
  wire [1-1:0] stream_conv2d_4_parameter_14_data;
  wire [16-1:0] stream_conv2d_4_source_15_data;
  wire [1-1:0] stream_conv2d_4_parameter_16_data;
  wire [1-1:0] stream_conv2d_4_parameter_17_data;
  wire [5-1:0] stream_conv2d_4_parameter_18_data;
  wire [1-1:0] stream_conv2d_4_parameter_19_data;
  wire [16-1:0] stream_conv2d_4_source_20_data;
  wire [16-1:0] stream_conv2d_4_source_21_data;
  wire [16-1:0] stream_conv2d_4_source_22_data;
  wire [16-1:0] stream_conv2d_4_source_23_data;
  wire [16-1:0] stream_conv2d_4_source_24_data;
  wire [16-1:0] stream_conv2d_4_source_25_data;
  wire [16-1:0] stream_conv2d_4_source_26_data;
  wire [16-1:0] stream_conv2d_4_source_27_data;
  wire [16-1:0] stream_conv2d_4_source_28_data;
  wire [16-1:0] stream_conv2d_4_source_29_data;
  wire [16-1:0] stream_conv2d_4_source_30_data;
  wire [16-1:0] stream_conv2d_4_source_31_data;
  wire [16-1:0] stream_conv2d_4_source_32_data;
  wire [16-1:0] stream_conv2d_4_source_33_data;
  wire [16-1:0] stream_conv2d_4_source_34_data;
  wire [16-1:0] stream_conv2d_4_source_35_data;
  wire [16-1:0] stream_conv2d_4_source_36_data;
  wire [16-1:0] stream_conv2d_4_source_37_data;
  reg __stream_conv2d_4_stream_ivalid_1;
  reg __stream_conv2d_4_stream_ivalid_2;
  reg __stream_conv2d_4_stream_ivalid_3;
  reg __stream_conv2d_4_stream_ivalid_4;
  reg __stream_conv2d_4_stream_ivalid_5;
  reg __stream_conv2d_4_stream_ivalid_6;
  reg __stream_conv2d_4_stream_ivalid_7;
  reg __stream_conv2d_4_stream_ivalid_8;
  reg __stream_conv2d_4_stream_ivalid_9;
  reg __stream_conv2d_4_stream_ivalid_10;
  reg __stream_conv2d_4_stream_ivalid_11;
  reg __stream_conv2d_4_stream_ivalid_12;
  reg __stream_conv2d_4_stream_ivalid_13;
  reg __stream_conv2d_4_stream_ivalid_14;
  reg __stream_conv2d_4_stream_ivalid_15;
  reg __stream_conv2d_4_stream_ivalid_16;
  reg __stream_conv2d_4_stream_ivalid_17;
  reg __stream_conv2d_4_stream_ivalid_18;
  reg __stream_conv2d_4_stream_ivalid_19;
  reg __stream_conv2d_4_stream_ivalid_20;
  reg __stream_conv2d_4_stream_ivalid_21;
  reg __stream_conv2d_4_stream_ivalid_22;
  reg __stream_conv2d_4_stream_ivalid_23;
  reg __stream_conv2d_4_stream_ivalid_24;
  reg __stream_conv2d_4_stream_ivalid_25;
  reg __stream_conv2d_4_stream_ivalid_26;
  reg __stream_conv2d_4_stream_ivalid_27;
  reg __stream_conv2d_4_stream_ivalid_28;
  reg __stream_conv2d_4_stream_ivalid_29;
  reg __stream_conv2d_4_stream_ivalid_30;
  reg __stream_conv2d_4_stream_ivalid_31;
  wire [16-1:0] _slice_data_1567;
  assign _slice_data_1567 = stream_conv2d_4_source_7_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_1568;
  assign _reinterpretcast_src_1568 = _slice_data_1567;
  wire signed [16-1:0] _reinterpretcast_data_1568;
  assign _reinterpretcast_data_1568 = _reinterpretcast_src_1568;
  wire signed [16-1:0] _cond_data_1569;
  assign _cond_data_1569 = (stream_conv2d_4_parameter_6_data)? _reinterpretcast_data_1568 : _reinterpretcast_data_1568;
  wire [16-1:0] _slice_data_1574;
  assign _slice_data_1574 = stream_conv2d_4_source_9_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_1575;
  assign _reinterpretcast_src_1575 = _slice_data_1574;
  wire signed [16-1:0] _reinterpretcast_data_1575;
  assign _reinterpretcast_data_1575 = _reinterpretcast_src_1575;
  wire signed [16-1:0] _cond_data_1576;
  assign _cond_data_1576 = (stream_conv2d_4_parameter_8_data)? _reinterpretcast_data_1575 : _reinterpretcast_data_1575;
  wire [16-1:0] _slice_data_1581;
  assign _slice_data_1581 = stream_conv2d_4_source_11_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_1582;
  assign _reinterpretcast_src_1582 = _slice_data_1581;
  wire [16-1:0] _reinterpretcast_data_1582;
  assign _reinterpretcast_data_1582 = _reinterpretcast_src_1582;
  wire [16-1:0] _cond_data_1583;
  assign _cond_data_1583 = (stream_conv2d_4_parameter_10_data)? _reinterpretcast_data_1582 : _reinterpretcast_data_1582;
  wire [16-1:0] _slice_data_1588;
  assign _slice_data_1588 = stream_conv2d_4_source_13_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_1589;
  assign _reinterpretcast_src_1589 = _slice_data_1588;
  wire [16-1:0] _reinterpretcast_data_1589;
  assign _reinterpretcast_data_1589 = _reinterpretcast_src_1589;
  wire [16-1:0] _cond_data_1590;
  assign _cond_data_1590 = (stream_conv2d_4_parameter_12_data)? _reinterpretcast_data_1589 : _reinterpretcast_data_1589;
  wire [16-1:0] _slice_data_1595;
  assign _slice_data_1595 = stream_conv2d_4_source_15_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_1596;
  assign _reinterpretcast_src_1596 = _slice_data_1595;
  wire [16-1:0] _reinterpretcast_data_1596;
  assign _reinterpretcast_data_1596 = _reinterpretcast_src_1596;
  wire [16-1:0] _cond_data_1597;
  assign _cond_data_1597 = (stream_conv2d_4_parameter_14_data)? _reinterpretcast_data_1596 : _reinterpretcast_data_1596;
  reg [1-1:0] _eq_data_1611;
  reg [1-1:0] _eq_data_1615;
  reg [1-1:0] _eq_data_1618;
  reg [1-1:0] _eq_data_1621;
  reg [1-1:0] _eq_data_1625;
  reg [1-1:0] _eq_data_1628;
  reg [1-1:0] _eq_data_1631;
  reg [1-1:0] _eq_data_1635;
  reg [1-1:0] _eq_data_1638;
  reg [1-1:0] _eq_data_1641;
  reg [1-1:0] _eq_data_1645;
  reg [1-1:0] _eq_data_1648;
  reg [1-1:0] _eq_data_1651;
  reg [1-1:0] _eq_data_1655;
  reg [1-1:0] _eq_data_1658;
  reg [1-1:0] _eq_data_1661;
  reg [1-1:0] _eq_data_1665;
  reg [1-1:0] _eq_data_1668;
  reg [1-1:0] _eq_data_1671;
  reg [1-1:0] _eq_data_1675;
  reg [1-1:0] _eq_data_1678;
  reg [1-1:0] _eq_data_1681;
  reg [1-1:0] _eq_data_1685;
  reg [1-1:0] _eq_data_1688;
  reg [1-1:0] _eq_data_1691;
  reg [1-1:0] _eq_data_1695;
  reg [1-1:0] _eq_data_1698;
  reg [1-1:0] _eq_data_1701;
  reg [1-1:0] _eq_data_1705;
  reg [1-1:0] _eq_data_1708;
  reg [1-1:0] _eq_data_1711;
  reg [1-1:0] _eq_data_1715;
  reg [1-1:0] _eq_data_1718;
  reg [1-1:0] _eq_data_1721;
  reg [1-1:0] _eq_data_1725;
  reg [1-1:0] _eq_data_1728;
  reg [1-1:0] _eq_data_1731;
  reg [1-1:0] _eq_data_1735;
  reg [1-1:0] _eq_data_1738;
  reg [1-1:0] _eq_data_1741;
  reg [1-1:0] _eq_data_1745;
  reg [1-1:0] _eq_data_1748;
  reg [1-1:0] _eq_data_1751;
  reg [1-1:0] _eq_data_1755;
  reg [1-1:0] _eq_data_1758;
  reg [1-1:0] _eq_data_1761;
  reg [1-1:0] _eq_data_1765;
  reg [1-1:0] _eq_data_1768;
  reg [1-1:0] _eq_data_1771;
  reg [1-1:0] _eq_data_1775;
  reg [1-1:0] _eq_data_1778;
  reg [1-1:0] _eq_data_1781;
  reg [1-1:0] _eq_data_1785;
  reg [1-1:0] _eq_data_1788;
  wire [16-1:0] _reinterpretcast_src_1881;
  assign _reinterpretcast_src_1881 = stream_conv2d_4_source_29_data;
  wire signed [16-1:0] _reinterpretcast_data_1881;
  assign _reinterpretcast_data_1881 = _reinterpretcast_src_1881;
  wire [16-1:0] _reinterpretcast_src_1882;
  assign _reinterpretcast_src_1882 = stream_conv2d_4_source_30_data;
  wire signed [16-1:0] _reinterpretcast_data_1882;
  assign _reinterpretcast_data_1882 = _reinterpretcast_src_1882;
  wire [16-1:0] _reinterpretcast_src_1883;
  assign _reinterpretcast_src_1883 = stream_conv2d_4_source_31_data;
  wire signed [16-1:0] _reinterpretcast_data_1883;
  assign _reinterpretcast_data_1883 = _reinterpretcast_src_1883;
  wire [16-1:0] _reinterpretcast_src_1884;
  assign _reinterpretcast_src_1884 = stream_conv2d_4_source_32_data;
  wire signed [16-1:0] _reinterpretcast_data_1884;
  assign _reinterpretcast_data_1884 = _reinterpretcast_src_1884;
  wire [16-1:0] _reinterpretcast_src_1885;
  assign _reinterpretcast_src_1885 = stream_conv2d_4_source_33_data;
  wire signed [16-1:0] _reinterpretcast_data_1885;
  assign _reinterpretcast_data_1885 = _reinterpretcast_src_1885;
  wire [16-1:0] _reinterpretcast_src_1886;
  assign _reinterpretcast_src_1886 = stream_conv2d_4_source_34_data;
  wire signed [16-1:0] _reinterpretcast_data_1886;
  assign _reinterpretcast_data_1886 = _reinterpretcast_src_1886;
  wire [16-1:0] _reinterpretcast_src_1887;
  assign _reinterpretcast_src_1887 = stream_conv2d_4_source_35_data;
  wire signed [16-1:0] _reinterpretcast_data_1887;
  assign _reinterpretcast_data_1887 = _reinterpretcast_src_1887;
  wire [16-1:0] _reinterpretcast_src_1888;
  assign _reinterpretcast_src_1888 = stream_conv2d_4_source_36_data;
  wire signed [16-1:0] _reinterpretcast_data_1888;
  assign _reinterpretcast_data_1888 = _reinterpretcast_src_1888;
  wire [16-1:0] _reinterpretcast_src_1889;
  assign _reinterpretcast_src_1889 = stream_conv2d_4_source_37_data;
  wire signed [16-1:0] _reinterpretcast_data_1889;
  assign _reinterpretcast_data_1889 = _reinterpretcast_src_1889;
  wire [1-1:0] _pointer_data_1890;
  assign _pointer_data_1890 = stream_conv2d_4_parameter_3_data[1'sd0];
  wire [1-1:0] _pointer_data_1892;
  assign _pointer_data_1892 = stream_conv2d_4_parameter_3_data[2'sd1];
  wire [1-1:0] _pointer_data_1894;
  assign _pointer_data_1894 = stream_conv2d_4_parameter_3_data[3'sd2];
  wire [1-1:0] _pointer_data_1896;
  assign _pointer_data_1896 = stream_conv2d_4_parameter_3_data[3'sd3];
  wire [1-1:0] _pointer_data_1898;
  assign _pointer_data_1898 = stream_conv2d_4_parameter_3_data[4'sd4];
  wire [1-1:0] _pointer_data_1900;
  assign _pointer_data_1900 = stream_conv2d_4_parameter_3_data[4'sd5];
  wire [1-1:0] _pointer_data_1902;
  assign _pointer_data_1902 = stream_conv2d_4_parameter_3_data[4'sd6];
  wire [1-1:0] _pointer_data_1904;
  assign _pointer_data_1904 = stream_conv2d_4_parameter_3_data[4'sd7];
  wire [1-1:0] _pointer_data_1906;
  assign _pointer_data_1906 = stream_conv2d_4_parameter_3_data[5'sd8];
  reg [16-1:0] _plus_data_1943;
  reg [16-1:0] _plus_data_1962;
  reg [16-1:0] _plus_data_1981;
  reg [16-1:0] _plus_data_2000;
  reg [16-1:0] _plus_data_2019;
  reg [16-1:0] _plus_data_2038;
  reg [16-1:0] _plus_data_2057;
  reg [16-1:0] _plus_data_2076;
  reg [16-1:0] _plus_data_2095;
  reg [16-1:0] _plus_data_2111;
  reg [16-1:0] _plus_data_2130;
  reg [16-1:0] __delay_data_2258__variable_1604;
  reg [16-1:0] __delay_data_2259__variable_1603;
  reg [16-1:0] __delay_data_2260__variable_1602;
  reg [16-1:0] __delay_data_2261__variable_1607;
  reg [16-1:0] __delay_data_2262__variable_1606;
  reg [16-1:0] __delay_data_2263__variable_1605;
  reg [16-1:0] __delay_data_2264__variable_1610;
  reg [16-1:0] __delay_data_2265__variable_1609;
  reg [16-1:0] __delay_data_2266__variable_1608;
  reg [1-1:0] __delay_data_2267_pointer_1890;
  reg signed [16-1:0] __delay_data_2268_reinterpretcast_1881;
  reg [1-1:0] __delay_data_2269_pointer_1892;
  reg signed [16-1:0] __delay_data_2270_reinterpretcast_1882;
  reg [1-1:0] __delay_data_2271_pointer_1894;
  reg signed [16-1:0] __delay_data_2272_reinterpretcast_1883;
  reg [1-1:0] __delay_data_2273_pointer_1896;
  reg signed [16-1:0] __delay_data_2274_reinterpretcast_1884;
  reg [1-1:0] __delay_data_2275_pointer_1898;
  reg signed [16-1:0] __delay_data_2276_reinterpretcast_1885;
  reg [1-1:0] __delay_data_2277_pointer_1900;
  reg signed [16-1:0] __delay_data_2278_reinterpretcast_1886;
  reg [1-1:0] __delay_data_2279_pointer_1902;
  reg signed [16-1:0] __delay_data_2280_reinterpretcast_1887;
  reg [1-1:0] __delay_data_2281_pointer_1904;
  reg signed [16-1:0] __delay_data_2282_reinterpretcast_1888;
  reg [1-1:0] __delay_data_2283_pointer_1906;
  reg signed [16-1:0] __delay_data_2284_reinterpretcast_1889;
  reg [1-1:0] __delay_data_2285__variable_1553;
  reg [1-1:0] __delay_data_2310__variable_1548;
  reg signed [16-1:0] __delay_data_2323_cond_1569;
  reg signed [16-1:0] __delay_data_2342_cond_1576;
  wire signed [16-1:0] _cond_data_1613;
  assign _cond_data_1613 = (_eq_data_1611)? __delay_data_2258__variable_1604 : 1'sd0;
  wire signed [16-1:0] _cond_data_1617;
  assign _cond_data_1617 = (_eq_data_1615)? __delay_data_2259__variable_1603 : _cond_data_1613;
  wire signed [16-1:0] _cond_data_1620;
  assign _cond_data_1620 = (_eq_data_1618)? __delay_data_2260__variable_1602 : _cond_data_1617;
  wire signed [16-1:0] _cond_data_1623;
  assign _cond_data_1623 = (_eq_data_1621)? __delay_data_2260__variable_1602 : 1'sd0;
  wire signed [16-1:0] _cond_data_1627;
  assign _cond_data_1627 = (_eq_data_1625)? __delay_data_2258__variable_1604 : _cond_data_1623;
  wire signed [16-1:0] _cond_data_1630;
  assign _cond_data_1630 = (_eq_data_1628)? __delay_data_2259__variable_1603 : _cond_data_1627;
  wire signed [16-1:0] _cond_data_1633;
  assign _cond_data_1633 = (_eq_data_1631)? __delay_data_2259__variable_1603 : 1'sd0;
  wire signed [16-1:0] _cond_data_1637;
  assign _cond_data_1637 = (_eq_data_1635)? __delay_data_2260__variable_1602 : _cond_data_1633;
  wire signed [16-1:0] _cond_data_1640;
  assign _cond_data_1640 = (_eq_data_1638)? __delay_data_2258__variable_1604 : _cond_data_1637;
  wire signed [16-1:0] _cond_data_1643;
  assign _cond_data_1643 = (_eq_data_1641)? __delay_data_2261__variable_1607 : 1'sd0;
  wire signed [16-1:0] _cond_data_1647;
  assign _cond_data_1647 = (_eq_data_1645)? __delay_data_2262__variable_1606 : _cond_data_1643;
  wire signed [16-1:0] _cond_data_1650;
  assign _cond_data_1650 = (_eq_data_1648)? __delay_data_2263__variable_1605 : _cond_data_1647;
  wire signed [16-1:0] _cond_data_1653;
  assign _cond_data_1653 = (_eq_data_1651)? __delay_data_2263__variable_1605 : 1'sd0;
  wire signed [16-1:0] _cond_data_1657;
  assign _cond_data_1657 = (_eq_data_1655)? __delay_data_2261__variable_1607 : _cond_data_1653;
  wire signed [16-1:0] _cond_data_1660;
  assign _cond_data_1660 = (_eq_data_1658)? __delay_data_2262__variable_1606 : _cond_data_1657;
  wire signed [16-1:0] _cond_data_1663;
  assign _cond_data_1663 = (_eq_data_1661)? __delay_data_2262__variable_1606 : 1'sd0;
  wire signed [16-1:0] _cond_data_1667;
  assign _cond_data_1667 = (_eq_data_1665)? __delay_data_2263__variable_1605 : _cond_data_1663;
  wire signed [16-1:0] _cond_data_1670;
  assign _cond_data_1670 = (_eq_data_1668)? __delay_data_2261__variable_1607 : _cond_data_1667;
  wire signed [16-1:0] _cond_data_1673;
  assign _cond_data_1673 = (_eq_data_1671)? __delay_data_2264__variable_1610 : 1'sd0;
  wire signed [16-1:0] _cond_data_1677;
  assign _cond_data_1677 = (_eq_data_1675)? __delay_data_2265__variable_1609 : _cond_data_1673;
  wire signed [16-1:0] _cond_data_1680;
  assign _cond_data_1680 = (_eq_data_1678)? __delay_data_2266__variable_1608 : _cond_data_1677;
  wire signed [16-1:0] _cond_data_1683;
  assign _cond_data_1683 = (_eq_data_1681)? __delay_data_2266__variable_1608 : 1'sd0;
  wire signed [16-1:0] _cond_data_1687;
  assign _cond_data_1687 = (_eq_data_1685)? __delay_data_2264__variable_1610 : _cond_data_1683;
  wire signed [16-1:0] _cond_data_1690;
  assign _cond_data_1690 = (_eq_data_1688)? __delay_data_2265__variable_1609 : _cond_data_1687;
  wire signed [16-1:0] _cond_data_1693;
  assign _cond_data_1693 = (_eq_data_1691)? __delay_data_2265__variable_1609 : 1'sd0;
  wire signed [16-1:0] _cond_data_1697;
  assign _cond_data_1697 = (_eq_data_1695)? __delay_data_2266__variable_1608 : _cond_data_1693;
  wire signed [16-1:0] _cond_data_1700;
  assign _cond_data_1700 = (_eq_data_1698)? __delay_data_2264__variable_1610 : _cond_data_1697;
  wire signed [16-1:0] _cond_data_1703;
  assign _cond_data_1703 = (_eq_data_1701)? _cond_data_1680 : 1'sd0;
  wire signed [16-1:0] _cond_data_1707;
  assign _cond_data_1707 = (_eq_data_1705)? _cond_data_1650 : _cond_data_1703;
  wire signed [16-1:0] _cond_data_1710;
  assign _cond_data_1710 = (_eq_data_1708)? _cond_data_1620 : _cond_data_1707;
  wire signed [16-1:0] _cond_data_1713;
  assign _cond_data_1713 = (_eq_data_1711)? _cond_data_1620 : 1'sd0;
  wire signed [16-1:0] _cond_data_1717;
  assign _cond_data_1717 = (_eq_data_1715)? _cond_data_1680 : _cond_data_1713;
  wire signed [16-1:0] _cond_data_1720;
  assign _cond_data_1720 = (_eq_data_1718)? _cond_data_1650 : _cond_data_1717;
  wire signed [16-1:0] _cond_data_1723;
  assign _cond_data_1723 = (_eq_data_1721)? _cond_data_1650 : 1'sd0;
  wire signed [16-1:0] _cond_data_1727;
  assign _cond_data_1727 = (_eq_data_1725)? _cond_data_1620 : _cond_data_1723;
  wire signed [16-1:0] _cond_data_1730;
  assign _cond_data_1730 = (_eq_data_1728)? _cond_data_1680 : _cond_data_1727;
  wire signed [16-1:0] _cond_data_1733;
  assign _cond_data_1733 = (_eq_data_1731)? _cond_data_1690 : 1'sd0;
  wire signed [16-1:0] _cond_data_1737;
  assign _cond_data_1737 = (_eq_data_1735)? _cond_data_1660 : _cond_data_1733;
  wire signed [16-1:0] _cond_data_1740;
  assign _cond_data_1740 = (_eq_data_1738)? _cond_data_1630 : _cond_data_1737;
  wire signed [16-1:0] _cond_data_1743;
  assign _cond_data_1743 = (_eq_data_1741)? _cond_data_1630 : 1'sd0;
  wire signed [16-1:0] _cond_data_1747;
  assign _cond_data_1747 = (_eq_data_1745)? _cond_data_1690 : _cond_data_1743;
  wire signed [16-1:0] _cond_data_1750;
  assign _cond_data_1750 = (_eq_data_1748)? _cond_data_1660 : _cond_data_1747;
  wire signed [16-1:0] _cond_data_1753;
  assign _cond_data_1753 = (_eq_data_1751)? _cond_data_1660 : 1'sd0;
  wire signed [16-1:0] _cond_data_1757;
  assign _cond_data_1757 = (_eq_data_1755)? _cond_data_1630 : _cond_data_1753;
  wire signed [16-1:0] _cond_data_1760;
  assign _cond_data_1760 = (_eq_data_1758)? _cond_data_1690 : _cond_data_1757;
  wire signed [16-1:0] _cond_data_1763;
  assign _cond_data_1763 = (_eq_data_1761)? _cond_data_1700 : 1'sd0;
  wire signed [16-1:0] _cond_data_1767;
  assign _cond_data_1767 = (_eq_data_1765)? _cond_data_1670 : _cond_data_1763;
  wire signed [16-1:0] _cond_data_1770;
  assign _cond_data_1770 = (_eq_data_1768)? _cond_data_1640 : _cond_data_1767;
  wire signed [16-1:0] _cond_data_1773;
  assign _cond_data_1773 = (_eq_data_1771)? _cond_data_1640 : 1'sd0;
  wire signed [16-1:0] _cond_data_1777;
  assign _cond_data_1777 = (_eq_data_1775)? _cond_data_1700 : _cond_data_1773;
  wire signed [16-1:0] _cond_data_1780;
  assign _cond_data_1780 = (_eq_data_1778)? _cond_data_1670 : _cond_data_1777;
  wire signed [16-1:0] _cond_data_1783;
  assign _cond_data_1783 = (_eq_data_1781)? _cond_data_1670 : 1'sd0;
  wire signed [16-1:0] _cond_data_1787;
  assign _cond_data_1787 = (_eq_data_1785)? _cond_data_1640 : _cond_data_1783;
  wire signed [16-1:0] _cond_data_1790;
  assign _cond_data_1790 = (_eq_data_1788)? _cond_data_1700 : _cond_data_1787;
  wire signed [16-1:0] _reinterpretcast_src_1827;
  assign _reinterpretcast_src_1827 = _cond_data_1710;
  wire signed [16-1:0] _reinterpretcast_data_1827;
  assign _reinterpretcast_data_1827 = _reinterpretcast_src_1827;
  wire signed [16-1:0] _reinterpretcast_src_1828;
  assign _reinterpretcast_src_1828 = _cond_data_1740;
  wire signed [16-1:0] _reinterpretcast_data_1828;
  assign _reinterpretcast_data_1828 = _reinterpretcast_src_1828;
  wire signed [16-1:0] _reinterpretcast_src_1829;
  assign _reinterpretcast_src_1829 = _cond_data_1770;
  wire signed [16-1:0] _reinterpretcast_data_1829;
  assign _reinterpretcast_data_1829 = _reinterpretcast_src_1829;
  wire signed [16-1:0] _reinterpretcast_src_1830;
  assign _reinterpretcast_src_1830 = _cond_data_1720;
  wire signed [16-1:0] _reinterpretcast_data_1830;
  assign _reinterpretcast_data_1830 = _reinterpretcast_src_1830;
  wire signed [16-1:0] _reinterpretcast_src_1831;
  assign _reinterpretcast_src_1831 = _cond_data_1750;
  wire signed [16-1:0] _reinterpretcast_data_1831;
  assign _reinterpretcast_data_1831 = _reinterpretcast_src_1831;
  wire signed [16-1:0] _reinterpretcast_src_1832;
  assign _reinterpretcast_src_1832 = _cond_data_1780;
  wire signed [16-1:0] _reinterpretcast_data_1832;
  assign _reinterpretcast_data_1832 = _reinterpretcast_src_1832;
  wire signed [16-1:0] _reinterpretcast_src_1833;
  assign _reinterpretcast_src_1833 = _cond_data_1730;
  wire signed [16-1:0] _reinterpretcast_data_1833;
  assign _reinterpretcast_data_1833 = _reinterpretcast_src_1833;
  wire signed [16-1:0] _reinterpretcast_src_1834;
  assign _reinterpretcast_src_1834 = _cond_data_1760;
  wire signed [16-1:0] _reinterpretcast_data_1834;
  assign _reinterpretcast_data_1834 = _reinterpretcast_src_1834;
  wire signed [16-1:0] _reinterpretcast_src_1835;
  assign _reinterpretcast_src_1835 = _cond_data_1790;
  wire signed [16-1:0] _reinterpretcast_data_1835;
  assign _reinterpretcast_data_1835 = _reinterpretcast_src_1835;
  wire signed [16-1:0] _cond_data_1909;
  assign _cond_data_1909 = (__delay_data_2267_pointer_1890)? 1'sd0 : _reinterpretcast_data_1827;
  wire signed [16-1:0] _cond_data_1911;
  assign _cond_data_1911 = (__delay_data_2269_pointer_1892)? 1'sd0 : _reinterpretcast_data_1828;
  wire signed [16-1:0] _cond_data_1913;
  assign _cond_data_1913 = (__delay_data_2271_pointer_1894)? 1'sd0 : _reinterpretcast_data_1829;
  wire signed [16-1:0] _cond_data_1915;
  assign _cond_data_1915 = (__delay_data_2273_pointer_1896)? 1'sd0 : _reinterpretcast_data_1830;
  wire signed [16-1:0] _cond_data_1917;
  assign _cond_data_1917 = (__delay_data_2275_pointer_1898)? 1'sd0 : _reinterpretcast_data_1831;
  wire signed [16-1:0] _cond_data_1919;
  assign _cond_data_1919 = (__delay_data_2277_pointer_1900)? 1'sd0 : _reinterpretcast_data_1832;
  wire signed [16-1:0] _cond_data_1921;
  assign _cond_data_1921 = (__delay_data_2279_pointer_1902)? 1'sd0 : _reinterpretcast_data_1833;
  wire signed [16-1:0] _cond_data_1923;
  assign _cond_data_1923 = (__delay_data_2281_pointer_1904)? 1'sd0 : _reinterpretcast_data_1834;
  wire signed [16-1:0] _cond_data_1925;
  assign _cond_data_1925 = (__delay_data_2283_pointer_1906)? 1'sd0 : _reinterpretcast_data_1835;
  reg signed [16-1:0] __variable_wdata_1352;
  assign mul_18_x_data = __variable_wdata_1352;
  reg signed [16-1:0] __variable_wdata_1353;
  assign mul_18_y_data = __variable_wdata_1353;
  reg [5-1:0] __variable_wdata_1354;
  assign mul_18_rshift_data = __variable_wdata_1354;
  reg signed [16-1:0] __variable_wdata_1373;
  assign mul_19_x_data = __variable_wdata_1373;
  reg signed [16-1:0] __variable_wdata_1374;
  assign mul_19_y_data = __variable_wdata_1374;
  reg [5-1:0] __variable_wdata_1375;
  assign mul_19_rshift_data = __variable_wdata_1375;
  assign _mul_19_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _mul_19_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_19_stream_internal_oready;
  reg signed [16-1:0] __variable_wdata_1394;
  assign mul_20_x_data = __variable_wdata_1394;
  reg signed [16-1:0] __variable_wdata_1395;
  assign mul_20_y_data = __variable_wdata_1395;
  reg [5-1:0] __variable_wdata_1396;
  assign mul_20_rshift_data = __variable_wdata_1396;
  assign _mul_20_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _mul_20_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_20_stream_internal_oready;
  reg signed [16-1:0] __variable_wdata_1415;
  assign mul_21_x_data = __variable_wdata_1415;
  reg signed [16-1:0] __variable_wdata_1416;
  assign mul_21_y_data = __variable_wdata_1416;
  reg [5-1:0] __variable_wdata_1417;
  assign mul_21_rshift_data = __variable_wdata_1417;
  assign _mul_21_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _mul_21_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_21_stream_internal_oready;
  reg signed [16-1:0] __variable_wdata_1436;
  assign mul_22_x_data = __variable_wdata_1436;
  reg signed [16-1:0] __variable_wdata_1437;
  assign mul_22_y_data = __variable_wdata_1437;
  reg [5-1:0] __variable_wdata_1438;
  assign mul_22_rshift_data = __variable_wdata_1438;
  assign _mul_22_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _mul_22_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_22_stream_internal_oready;
  reg signed [16-1:0] __variable_wdata_1457;
  assign mul_23_x_data = __variable_wdata_1457;
  reg signed [16-1:0] __variable_wdata_1458;
  assign mul_23_y_data = __variable_wdata_1458;
  reg [5-1:0] __variable_wdata_1459;
  assign mul_23_rshift_data = __variable_wdata_1459;
  assign _mul_23_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _mul_23_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_23_stream_internal_oready;
  reg signed [16-1:0] __variable_wdata_1478;
  assign mul_24_x_data = __variable_wdata_1478;
  reg signed [16-1:0] __variable_wdata_1479;
  assign mul_24_y_data = __variable_wdata_1479;
  reg [5-1:0] __variable_wdata_1480;
  assign mul_24_rshift_data = __variable_wdata_1480;
  assign _mul_24_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _mul_24_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_24_stream_internal_oready;
  reg signed [16-1:0] __variable_wdata_1499;
  assign mul_25_x_data = __variable_wdata_1499;
  reg signed [16-1:0] __variable_wdata_1500;
  assign mul_25_y_data = __variable_wdata_1500;
  reg [5-1:0] __variable_wdata_1501;
  assign mul_25_rshift_data = __variable_wdata_1501;
  assign _mul_25_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _mul_25_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_25_stream_internal_oready;
  reg signed [16-1:0] __variable_wdata_1520;
  assign mul_26_x_data = __variable_wdata_1520;
  reg signed [16-1:0] __variable_wdata_1521;
  assign mul_26_y_data = __variable_wdata_1521;
  reg [5-1:0] __variable_wdata_1522;
  assign mul_26_rshift_data = __variable_wdata_1522;
  assign _mul_26_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _mul_26_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_26_stream_internal_oready;
  reg [1-1:0] __delay_data_2286__delay_2285__variable_1553;
  reg [16-1:0] __delay_data_2298_plus_2111;
  reg [1-1:0] __delay_data_2311__delay_2310__variable_1548;
  reg signed [16-1:0] __delay_data_2324__delay_2323_cond_1569;
  reg signed [16-1:0] __delay_data_2343__delay_2342_cond_1576;
  reg [16-1:0] __delay_data_2362_plus_2130;
  reg [1-1:0] __delay_data_2287__delay_2286__delay_2285__variable_1553;
  reg [16-1:0] __delay_data_2299__delay_2298_plus_2111;
  reg [1-1:0] __delay_data_2312__delay_2311__delay_2310__variable_1548;
  reg signed [16-1:0] __delay_data_2325__delay_2324__delay_2323_cond_1569;
  reg signed [16-1:0] __delay_data_2344__delay_2343__delay_2342_cond_1576;
  reg [16-1:0] __delay_data_2363__delay_2362_plus_2130;
  reg [1-1:0] __delay_data_2288__delay_2287__delay_2286____variable_1553;
  reg [16-1:0] __delay_data_2300__delay_2299__delay_2298_plus_2111;
  reg [1-1:0] __delay_data_2313__delay_2312__delay_2311____variable_1548;
  reg signed [16-1:0] __delay_data_2326__delay_2325__delay_2324___cond_1569;
  reg signed [16-1:0] __delay_data_2345__delay_2344__delay_2343___cond_1576;
  reg [16-1:0] __delay_data_2364__delay_2363__delay_2362_plus_2130;
  reg [1-1:0] __delay_data_2289__delay_2288__delay_2287____variable_1553;
  reg [16-1:0] __delay_data_2301__delay_2300__delay_2299___plus_2111;
  reg [1-1:0] __delay_data_2314__delay_2313__delay_2312____variable_1548;
  reg signed [16-1:0] __delay_data_2327__delay_2326__delay_2325___cond_1569;
  reg signed [16-1:0] __delay_data_2346__delay_2345__delay_2344___cond_1576;
  reg [16-1:0] __delay_data_2365__delay_2364__delay_2363___plus_2130;
  reg [1-1:0] __delay_data_2290__delay_2289__delay_2288____variable_1553;
  reg [16-1:0] __delay_data_2302__delay_2301__delay_2300___plus_2111;
  reg [1-1:0] __delay_data_2315__delay_2314__delay_2313____variable_1548;
  reg signed [16-1:0] __delay_data_2328__delay_2327__delay_2326___cond_1569;
  reg signed [16-1:0] __delay_data_2347__delay_2346__delay_2345___cond_1576;
  reg [16-1:0] __delay_data_2366__delay_2365__delay_2364___plus_2130;
  reg [1-1:0] __delay_data_2291__delay_2290__delay_2289____variable_1553;
  reg [16-1:0] __delay_data_2303__delay_2302__delay_2301___plus_2111;
  reg [1-1:0] __delay_data_2316__delay_2315__delay_2314____variable_1548;
  reg signed [16-1:0] __delay_data_2329__delay_2328__delay_2327___cond_1569;
  reg signed [16-1:0] __delay_data_2348__delay_2347__delay_2346___cond_1576;
  reg [16-1:0] __delay_data_2367__delay_2366__delay_2365___plus_2130;
  reg [1-1:0] __delay_data_2292__delay_2291__delay_2290____variable_1553;
  reg [16-1:0] __delay_data_2304__delay_2303__delay_2302___plus_2111;
  reg [1-1:0] __delay_data_2317__delay_2316__delay_2315____variable_1548;
  reg signed [16-1:0] __delay_data_2330__delay_2329__delay_2328___cond_1569;
  reg signed [16-1:0] __delay_data_2349__delay_2348__delay_2347___cond_1576;
  reg [16-1:0] __delay_data_2368__delay_2367__delay_2366___plus_2130;
  reg [1-1:0] __delay_data_2293__delay_2292__delay_2291____variable_1553;
  reg [16-1:0] __delay_data_2305__delay_2304__delay_2303___plus_2111;
  reg [1-1:0] __delay_data_2318__delay_2317__delay_2316____variable_1548;
  reg signed [16-1:0] __delay_data_2331__delay_2330__delay_2329___cond_1569;
  reg signed [16-1:0] __delay_data_2350__delay_2349__delay_2348___cond_1576;
  reg [16-1:0] __delay_data_2369__delay_2368__delay_2367___plus_2130;
  reg [1-1:0] __delay_data_2294__delay_2293__delay_2292____variable_1553;
  reg [16-1:0] __delay_data_2306__delay_2305__delay_2304___plus_2111;
  reg [1-1:0] __delay_data_2319__delay_2318__delay_2317____variable_1548;
  reg signed [16-1:0] __delay_data_2332__delay_2331__delay_2330___cond_1569;
  reg signed [16-1:0] __delay_data_2351__delay_2350__delay_2349___cond_1576;
  reg [16-1:0] __delay_data_2370__delay_2369__delay_2368___plus_2130;
  wire signed [32-1:0] __substreamoutput_data_1944;
  assign __substreamoutput_data_1944 = mul_18_z_data;
  wire signed [32-1:0] __substreamoutput_data_1963;
  assign __substreamoutput_data_1963 = mul_19_z_data;
  wire signed [32-1:0] __substreamoutput_data_1982;
  assign __substreamoutput_data_1982 = mul_20_z_data;
  wire signed [32-1:0] __substreamoutput_data_2001;
  assign __substreamoutput_data_2001 = mul_21_z_data;
  wire signed [32-1:0] __substreamoutput_data_2020;
  assign __substreamoutput_data_2020 = mul_22_z_data;
  wire signed [32-1:0] __substreamoutput_data_2039;
  assign __substreamoutput_data_2039 = mul_23_z_data;
  wire signed [32-1:0] __substreamoutput_data_2058;
  assign __substreamoutput_data_2058 = mul_24_z_data;
  wire signed [32-1:0] __substreamoutput_data_2077;
  assign __substreamoutput_data_2077 = mul_25_z_data;
  wire signed [32-1:0] __substreamoutput_data_2096;
  assign __substreamoutput_data_2096 = mul_26_z_data;
  reg signed [64-1:0] __variable_wdata_1304;
  assign add_tree_16_var0_data = __variable_wdata_1304;
  reg signed [64-1:0] __variable_wdata_1305;
  assign add_tree_16_var1_data = __variable_wdata_1305;
  reg signed [64-1:0] __variable_wdata_1306;
  assign add_tree_16_var2_data = __variable_wdata_1306;
  reg signed [64-1:0] __variable_wdata_1307;
  assign add_tree_16_var3_data = __variable_wdata_1307;
  reg signed [64-1:0] __variable_wdata_1308;
  assign add_tree_16_var4_data = __variable_wdata_1308;
  reg signed [64-1:0] __variable_wdata_1309;
  assign add_tree_16_var5_data = __variable_wdata_1309;
  reg signed [64-1:0] __variable_wdata_1310;
  assign add_tree_16_var6_data = __variable_wdata_1310;
  reg signed [64-1:0] __variable_wdata_1311;
  assign add_tree_16_var7_data = __variable_wdata_1311;
  reg signed [64-1:0] __variable_wdata_1312;
  assign add_tree_16_var8_data = __variable_wdata_1312;
  assign _add_tree_16_is_root = ((_stream_conv2d_4_busy)? 0 : 1) && 1;
  assign _add_tree_16_stream_oready = ((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _add_tree_16_stream_internal_oready;
  reg [1-1:0] __delay_data_2295__delay_2294__delay_2293____variable_1553;
  reg [16-1:0] __delay_data_2307__delay_2306__delay_2305___plus_2111;
  reg [1-1:0] __delay_data_2320__delay_2319__delay_2318____variable_1548;
  reg signed [16-1:0] __delay_data_2333__delay_2332__delay_2331___cond_1569;
  reg signed [16-1:0] __delay_data_2352__delay_2351__delay_2350___cond_1576;
  reg [16-1:0] __delay_data_2371__delay_2370__delay_2369___plus_2130;
  reg [1-1:0] __delay_data_2296__delay_2295__delay_2294____variable_1553;
  reg [16-1:0] __delay_data_2308__delay_2307__delay_2306___plus_2111;
  reg [1-1:0] __delay_data_2321__delay_2320__delay_2319____variable_1548;
  reg signed [16-1:0] __delay_data_2334__delay_2333__delay_2332___cond_1569;
  reg signed [16-1:0] __delay_data_2353__delay_2352__delay_2351___cond_1576;
  reg [16-1:0] __delay_data_2372__delay_2371__delay_2370___plus_2130;
  reg [1-1:0] __delay_data_2297__delay_2296__delay_2295____variable_1553;
  reg [16-1:0] __delay_data_2309__delay_2308__delay_2307___plus_2111;
  reg [1-1:0] __delay_data_2322__delay_2321__delay_2320____variable_1548;
  reg signed [16-1:0] __delay_data_2335__delay_2334__delay_2333___cond_1569;
  reg signed [16-1:0] __delay_data_2354__delay_2353__delay_2352___cond_1576;
  reg [16-1:0] __delay_data_2373__delay_2372__delay_2371___plus_2130;
  wire signed [64-1:0] __substreamoutput_data_2098;
  assign __substreamoutput_data_2098 = add_tree_16_sum_data;
  reg [1-1:0] __variable_wdata_1295;
  assign acc_14__reduce_reset_data = __variable_wdata_1295;
  reg signed [64-1:0] __variable_wdata_1280;
  assign acc_14_x_data = __variable_wdata_1280;
  reg [7-1:0] __variable_wdata_1281;
  assign acc_14_rshift_data = __variable_wdata_1281;
  reg [32-1:0] __variable_wdata_1282;
  assign acc_14_size_data = __variable_wdata_1282;
  reg signed [16-1:0] __delay_data_2336__delay_2335__delay_2334___cond_1569;
  reg signed [16-1:0] __delay_data_2355__delay_2354__delay_2353___cond_1576;
  reg [16-1:0] __delay_data_2374__delay_2373__delay_2372___plus_2130;
  reg signed [16-1:0] __delay_data_2337__delay_2336__delay_2335___cond_1569;
  reg signed [16-1:0] __delay_data_2356__delay_2355__delay_2354___cond_1576;
  reg [16-1:0] __delay_data_2375__delay_2374__delay_2373___plus_2130;
  reg signed [16-1:0] __delay_data_2338__delay_2337__delay_2336___cond_1569;
  reg signed [16-1:0] __delay_data_2357__delay_2356__delay_2355___cond_1576;
  reg [16-1:0] __delay_data_2376__delay_2375__delay_2374___plus_2130;
  reg signed [16-1:0] __delay_data_2339__delay_2338__delay_2337___cond_1569;
  reg signed [16-1:0] __delay_data_2358__delay_2357__delay_2356___cond_1576;
  reg [16-1:0] __delay_data_2377__delay_2376__delay_2375___plus_2130;
  reg signed [16-1:0] __delay_data_2340__delay_2339__delay_2338___cond_1569;
  reg signed [16-1:0] __delay_data_2359__delay_2358__delay_2357___cond_1576;
  reg [16-1:0] __delay_data_2378__delay_2377__delay_2376___plus_2130;
  reg signed [16-1:0] __delay_data_2341__delay_2340__delay_2339___cond_1569;
  reg signed [16-1:0] __delay_data_2360__delay_2359__delay_2358___cond_1576;
  reg [16-1:0] __delay_data_2379__delay_2378__delay_2377___plus_2130;
  wire signed [64-1:0] __substreamoutput_data_2112;
  assign __substreamoutput_data_2112 = acc_14_sum_data;
  wire [1-1:0] __substreamoutput_data_2113;
  assign __substreamoutput_data_2113 = acc_14_valid_data;
  reg signed [64-1:0] _plus_data_2114;
  reg signed [16-1:0] __delay_data_2361__delay_2360__delay_2359___cond_1576;
  reg [16-1:0] __delay_data_2380__delay_2379__delay_2378___plus_2130;
  reg [1-1:0] __delay_data_2382__substreamoutput_2113;
  reg signed [64-1:0] __variable_wdata_1318;
  assign mul_rshift_round_clip_17_x_data = __variable_wdata_1318;
  reg signed [16-1:0] __variable_wdata_1319;
  assign mul_rshift_round_clip_17_y_data = __variable_wdata_1319;
  reg [7-1:0] __variable_wdata_1320;
  assign mul_rshift_round_clip_17_rshift_data = __variable_wdata_1320;
  assign _stream_conv2d_4_stream_internal_oready = ((_stream_conv2d_4_busy)? _mul_rshift_round_clip_17_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _acc_14_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _add_tree_16_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_26_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_25_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_24_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_23_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_22_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_21_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_20_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_19_stream_internal_oready : 1) && (((_stream_conv2d_4_busy)? _mul_18_stream_internal_oready : 1) && 1)))))))))));
  reg [1-1:0] __delay_data_2383__delay_2382__substreamoutput_2113;
  reg [1-1:0] __delay_data_2384__delay_2383____substreamoutput_2113;
  reg [1-1:0] __delay_data_2385__delay_2384____substreamoutput_2113;
  reg [1-1:0] __delay_data_2386__delay_2385____substreamoutput_2113;
  reg [1-1:0] __delay_data_2387__delay_2386____substreamoutput_2113;
  reg [1-1:0] __delay_data_2388__delay_2387____substreamoutput_2113;
  reg [1-1:0] __delay_data_2389__delay_2388____substreamoutput_2113;
  reg [1-1:0] __delay_data_2390__delay_2389____substreamoutput_2113;
  reg [1-1:0] __delay_data_2391__delay_2390____substreamoutput_2113;
  wire signed [16-1:0] __substreamoutput_data_2131;
  assign __substreamoutput_data_2131 = mul_rshift_round_clip_17_z_data;
  reg [1-1:0] _greaterthan_data_2133;
  reg signed [16-1:0] __delay_data_2381__substreamoutput_2131;
  reg [1-1:0] __delay_data_2392__delay_2391____substreamoutput_2113;
  reg signed [16-1:0] _cond_data_2135;
  reg [1-1:0] __delay_data_2393__delay_2392____substreamoutput_2113;
  wire signed [16-1:0] _reinterpretcast_src_2136;
  assign _reinterpretcast_src_2136 = _cond_data_2135;
  wire signed [16-1:0] _reinterpretcast_data_2136;
  assign _reinterpretcast_data_2136 = _reinterpretcast_src_2136;
  wire signed [16-1:0] stream_conv2d_4_sink_50_data;
  assign stream_conv2d_4_sink_50_data = _reinterpretcast_data_2136;
  wire [1-1:0] stream_conv2d_4_sink_51_data;
  assign stream_conv2d_4_sink_51_data = __delay_data_2393__delay_2392____substreamoutput_2113;
  wire _set_flag_328;
  assign _set_flag_328 = conv2d_4_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_1548;
  assign stream_conv2d_4_parameter_0_data = __variable_wdata_1548;
  wire _set_flag_329;
  assign _set_flag_329 = conv2d_4_comp_fsm == 3;
  reg [2-1:0] __variable_wdata_1549;
  assign stream_conv2d_4_parameter_1_data = __variable_wdata_1549;
  wire _set_flag_330;
  assign _set_flag_330 = conv2d_4_comp_fsm == 3;
  reg [2-1:0] __variable_wdata_1550;
  assign stream_conv2d_4_parameter_2_data = __variable_wdata_1550;
  wire _set_flag_331;
  assign _set_flag_331 = conv2d_4_comp_fsm == 3;
  reg [9-1:0] __variable_wdata_1551;
  assign stream_conv2d_4_parameter_3_data = __variable_wdata_1551;
  wire _set_flag_332;
  assign _set_flag_332 = conv2d_4_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_1552;
  assign stream_conv2d_4_parameter_4_data = __variable_wdata_1552;
  wire _set_flag_333;
  assign _set_flag_333 = conv2d_4_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_1563;
  assign stream_conv2d_4_parameter_6_data = __variable_wdata_1563;
  reg [32-1:0] _source_stream_conv2d_4_source_7_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_7_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_7_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_7_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_7_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_7_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_7_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_7_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_7_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_7_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_7_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_7_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_7_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_7_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_7_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_7_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_7_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_7_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_7_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_7_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_7_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_7_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_7_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_7_pat_stride_buf_3;
  wire _set_flag_334;
  assign _set_flag_334 = conv2d_4_comp_fsm == 3;
  wire [1-1:0] read_rtl_bank_335;
  assign read_rtl_bank_335 = _stream_conv2d_4_source_7_source_ram_raddr;
  reg [1-1:0] _tmp_336;
  assign ram_w16_l512_id9_0_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_7_source_ram_renable && (_stream_conv2d_4_source_7_source_sel == 1))? _stream_conv2d_4_source_7_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id9_0_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_7_source_ram_renable && (_stream_conv2d_4_source_7_source_sel == 1))? 1'd1 : 0;
  localparam _tmp_337 = 1;
  wire [_tmp_337-1:0] _tmp_338;
  assign _tmp_338 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_7_source_ram_renable && (_stream_conv2d_4_source_7_source_sel == 1);
  reg [_tmp_337-1:0] __tmp_338_1;
  assign ram_w16_l512_id9_1_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_7_source_ram_renable && (_stream_conv2d_4_source_7_source_sel == 1))? _stream_conv2d_4_source_7_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id9_1_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_7_source_ram_renable && (_stream_conv2d_4_source_7_source_sel == 1))? 1'd1 : 0;
  localparam _tmp_339 = 1;
  wire [_tmp_339-1:0] _tmp_340;
  assign _tmp_340 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_7_source_ram_renable && (_stream_conv2d_4_source_7_source_sel == 1);
  reg [_tmp_339-1:0] __tmp_340_1;
  wire signed [16-1:0] read_rtl_rdata_341;
  wire read_rtl_rvalid_342;
  assign read_rtl_rdata_341 = (_tmp_336 == 0)? ram_w16_l512_id9_0_0_rdata : 
                              (_tmp_336 == 1)? ram_w16_l512_id9_1_0_rdata : 0;
  assign read_rtl_rvalid_342 = __tmp_338_1;
  assign _stream_conv2d_4_source_7_source_ram_rdata = (_stream_conv2d_4_source_7_source_sel == 1)? read_rtl_rdata_341 : 'hx;
  reg [16-1:0] __variable_wdata_1564;
  assign stream_conv2d_4_source_7_data = __variable_wdata_1564;
  reg [32-1:0] _stream_conv2d_4_source_7_source_pat_fsm_0;
  localparam _stream_conv2d_4_source_7_source_pat_fsm_0_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_7_source_pat_all_offset;
  assign _stream_conv2d_4_source_7_source_pat_all_offset = _stream_conv2d_4_source_7_source_offset_buf + _source_stream_conv2d_4_source_7_pat_cur_offset_0 + _source_stream_conv2d_4_source_7_pat_cur_offset_1 + _source_stream_conv2d_4_source_7_pat_cur_offset_2 + _source_stream_conv2d_4_source_7_pat_cur_offset_3;
  wire _set_flag_343;
  assign _set_flag_343 = conv2d_4_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_1570;
  assign stream_conv2d_4_parameter_8_data = __variable_wdata_1570;
  reg [32-1:0] _source_stream_conv2d_4_source_9_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_9_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_9_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_9_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_9_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_9_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_9_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_9_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_9_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_9_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_9_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_9_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_9_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_9_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_9_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_9_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_9_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_9_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_9_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_9_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_9_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_9_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_9_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_9_pat_stride_buf_3;
  wire _set_flag_344;
  assign _set_flag_344 = conv2d_4_comp_fsm == 3;
  wire [1-1:0] read_rtl_bank_345;
  assign read_rtl_bank_345 = _stream_conv2d_4_source_9_source_ram_raddr;
  reg [1-1:0] _tmp_346;
  assign ram_w16_l512_id10_0_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_9_source_ram_renable && (_stream_conv2d_4_source_9_source_sel == 2))? _stream_conv2d_4_source_9_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id10_0_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_9_source_ram_renable && (_stream_conv2d_4_source_9_source_sel == 2))? 1'd1 : 0;
  localparam _tmp_347 = 1;
  wire [_tmp_347-1:0] _tmp_348;
  assign _tmp_348 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_9_source_ram_renable && (_stream_conv2d_4_source_9_source_sel == 2);
  reg [_tmp_347-1:0] __tmp_348_1;
  assign ram_w16_l512_id10_1_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_9_source_ram_renable && (_stream_conv2d_4_source_9_source_sel == 2))? _stream_conv2d_4_source_9_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id10_1_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_9_source_ram_renable && (_stream_conv2d_4_source_9_source_sel == 2))? 1'd1 : 0;
  localparam _tmp_349 = 1;
  wire [_tmp_349-1:0] _tmp_350;
  assign _tmp_350 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_9_source_ram_renable && (_stream_conv2d_4_source_9_source_sel == 2);
  reg [_tmp_349-1:0] __tmp_350_1;
  wire signed [16-1:0] read_rtl_rdata_351;
  wire read_rtl_rvalid_352;
  assign read_rtl_rdata_351 = (_tmp_346 == 0)? ram_w16_l512_id10_0_0_rdata : 
                              (_tmp_346 == 1)? ram_w16_l512_id10_1_0_rdata : 0;
  assign read_rtl_rvalid_352 = __tmp_348_1;
  assign _stream_conv2d_4_source_9_source_ram_rdata = (_stream_conv2d_4_source_9_source_sel == 2)? read_rtl_rdata_351 : 'hx;
  reg [16-1:0] __variable_wdata_1571;
  assign stream_conv2d_4_source_9_data = __variable_wdata_1571;
  reg [32-1:0] _stream_conv2d_4_source_9_source_pat_fsm_1;
  localparam _stream_conv2d_4_source_9_source_pat_fsm_1_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_9_source_pat_all_offset;
  assign _stream_conv2d_4_source_9_source_pat_all_offset = _stream_conv2d_4_source_9_source_offset_buf + _source_stream_conv2d_4_source_9_pat_cur_offset_0 + _source_stream_conv2d_4_source_9_pat_cur_offset_1 + _source_stream_conv2d_4_source_9_pat_cur_offset_2 + _source_stream_conv2d_4_source_9_pat_cur_offset_3;
  wire _set_flag_353;
  assign _set_flag_353 = conv2d_4_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_1577;
  assign stream_conv2d_4_parameter_10_data = __variable_wdata_1577;
  wire _set_flag_354;
  assign _set_flag_354 = conv2d_4_comp_fsm == 3;
  reg [16-1:0] __variable_wdata_1578;
  assign stream_conv2d_4_source_11_data = __variable_wdata_1578;
  wire _set_flag_355;
  assign _set_flag_355 = conv2d_4_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_1584;
  assign stream_conv2d_4_parameter_12_data = __variable_wdata_1584;
  wire _set_flag_356;
  assign _set_flag_356 = conv2d_4_comp_fsm == 3;
  reg [16-1:0] __variable_wdata_1585;
  assign stream_conv2d_4_source_13_data = __variable_wdata_1585;
  wire _set_flag_357;
  assign _set_flag_357 = conv2d_4_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_1591;
  assign stream_conv2d_4_parameter_14_data = __variable_wdata_1591;
  wire _set_flag_358;
  assign _set_flag_358 = conv2d_4_comp_fsm == 3;
  reg [16-1:0] __variable_wdata_1592;
  assign stream_conv2d_4_source_15_data = __variable_wdata_1592;
  wire _set_flag_359;
  assign _set_flag_359 = conv2d_4_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_1598;
  assign stream_conv2d_4_parameter_16_data = __variable_wdata_1598;
  wire _set_flag_360;
  assign _set_flag_360 = conv2d_4_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_1599;
  assign stream_conv2d_4_parameter_17_data = __variable_wdata_1599;
  wire _set_flag_361;
  assign _set_flag_361 = conv2d_4_comp_fsm == 3;
  reg [5-1:0] __variable_wdata_1600;
  assign stream_conv2d_4_parameter_18_data = __variable_wdata_1600;
  wire _set_flag_362;
  assign _set_flag_362 = conv2d_4_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_1601;
  assign stream_conv2d_4_parameter_19_data = __variable_wdata_1601;
  reg [32-1:0] _source_stream_conv2d_4_source_20_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_20_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_20_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_20_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_20_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_20_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_20_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_20_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_20_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_20_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_20_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_20_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_20_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_20_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_20_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_20_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_20_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_20_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_20_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_20_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_20_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_20_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_20_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_20_pat_stride_buf_3;
  wire _set_flag_363;
  assign _set_flag_363 = conv2d_4_comp_fsm == 3;
  wire [1-1:0] read_rtl_bank_364;
  assign read_rtl_bank_364 = _stream_conv2d_4_source_20_source_ram_raddr;
  reg [1-1:0] _tmp_365;
  assign ram_w16_l512_id11_0_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_20_source_ram_renable && (_stream_conv2d_4_source_20_source_sel == 3))? _stream_conv2d_4_source_20_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id11_0_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_20_source_ram_renable && (_stream_conv2d_4_source_20_source_sel == 3))? 1'd1 : 0;
  localparam _tmp_366 = 1;
  wire [_tmp_366-1:0] _tmp_367;
  assign _tmp_367 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_20_source_ram_renable && (_stream_conv2d_4_source_20_source_sel == 3);
  reg [_tmp_366-1:0] __tmp_367_1;
  assign ram_w16_l512_id11_1_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_20_source_ram_renable && (_stream_conv2d_4_source_20_source_sel == 3))? _stream_conv2d_4_source_20_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id11_1_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_20_source_ram_renable && (_stream_conv2d_4_source_20_source_sel == 3))? 1'd1 : 0;
  localparam _tmp_368 = 1;
  wire [_tmp_368-1:0] _tmp_369;
  assign _tmp_369 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_20_source_ram_renable && (_stream_conv2d_4_source_20_source_sel == 3);
  reg [_tmp_368-1:0] __tmp_369_1;
  wire signed [16-1:0] read_rtl_rdata_370;
  wire read_rtl_rvalid_371;
  assign read_rtl_rdata_370 = (_tmp_365 == 0)? ram_w16_l512_id11_0_0_rdata : 
                              (_tmp_365 == 1)? ram_w16_l512_id11_1_0_rdata : 0;
  assign read_rtl_rvalid_371 = __tmp_367_1;
  assign _stream_conv2d_4_source_20_source_ram_rdata = (_stream_conv2d_4_source_20_source_sel == 3)? read_rtl_rdata_370 : 'hx;
  reg [16-1:0] __variable_wdata_1602;
  assign stream_conv2d_4_source_20_data = __variable_wdata_1602;
  reg [32-1:0] _stream_conv2d_4_source_20_source_pat_fsm_2;
  localparam _stream_conv2d_4_source_20_source_pat_fsm_2_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_20_source_pat_all_offset;
  assign _stream_conv2d_4_source_20_source_pat_all_offset = _stream_conv2d_4_source_20_source_offset_buf + _source_stream_conv2d_4_source_20_pat_cur_offset_0 + _source_stream_conv2d_4_source_20_pat_cur_offset_1 + _source_stream_conv2d_4_source_20_pat_cur_offset_2 + _source_stream_conv2d_4_source_20_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_21_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_21_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_21_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_21_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_21_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_21_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_21_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_21_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_21_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_21_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_21_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_21_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_21_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_21_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_21_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_21_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_21_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_21_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_21_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_21_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_21_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_21_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_21_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_21_pat_stride_buf_3;
  wire _set_flag_372;
  assign _set_flag_372 = conv2d_4_comp_fsm == 3;
  wire [1-1:0] read_rtl_bank_373;
  assign read_rtl_bank_373 = _stream_conv2d_4_source_21_source_ram_raddr;
  reg [1-1:0] _tmp_374;
  assign ram_w16_l512_id12_0_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_21_source_ram_renable && (_stream_conv2d_4_source_21_source_sel == 4))? _stream_conv2d_4_source_21_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id12_0_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_21_source_ram_renable && (_stream_conv2d_4_source_21_source_sel == 4))? 1'd1 : 0;
  localparam _tmp_375 = 1;
  wire [_tmp_375-1:0] _tmp_376;
  assign _tmp_376 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_21_source_ram_renable && (_stream_conv2d_4_source_21_source_sel == 4);
  reg [_tmp_375-1:0] __tmp_376_1;
  assign ram_w16_l512_id12_1_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_21_source_ram_renable && (_stream_conv2d_4_source_21_source_sel == 4))? _stream_conv2d_4_source_21_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id12_1_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_21_source_ram_renable && (_stream_conv2d_4_source_21_source_sel == 4))? 1'd1 : 0;
  localparam _tmp_377 = 1;
  wire [_tmp_377-1:0] _tmp_378;
  assign _tmp_378 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_21_source_ram_renable && (_stream_conv2d_4_source_21_source_sel == 4);
  reg [_tmp_377-1:0] __tmp_378_1;
  wire signed [16-1:0] read_rtl_rdata_379;
  wire read_rtl_rvalid_380;
  assign read_rtl_rdata_379 = (_tmp_374 == 0)? ram_w16_l512_id12_0_0_rdata : 
                              (_tmp_374 == 1)? ram_w16_l512_id12_1_0_rdata : 0;
  assign read_rtl_rvalid_380 = __tmp_376_1;
  assign _stream_conv2d_4_source_21_source_ram_rdata = (_stream_conv2d_4_source_21_source_sel == 4)? read_rtl_rdata_379 : 'hx;
  reg [16-1:0] __variable_wdata_1603;
  assign stream_conv2d_4_source_21_data = __variable_wdata_1603;
  reg [32-1:0] _stream_conv2d_4_source_21_source_pat_fsm_3;
  localparam _stream_conv2d_4_source_21_source_pat_fsm_3_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_21_source_pat_all_offset;
  assign _stream_conv2d_4_source_21_source_pat_all_offset = _stream_conv2d_4_source_21_source_offset_buf + _source_stream_conv2d_4_source_21_pat_cur_offset_0 + _source_stream_conv2d_4_source_21_pat_cur_offset_1 + _source_stream_conv2d_4_source_21_pat_cur_offset_2 + _source_stream_conv2d_4_source_21_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_22_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_22_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_22_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_22_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_22_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_22_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_22_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_22_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_22_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_22_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_22_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_22_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_22_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_22_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_22_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_22_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_22_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_22_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_22_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_22_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_22_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_22_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_22_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_22_pat_stride_buf_3;
  wire _set_flag_381;
  assign _set_flag_381 = conv2d_4_comp_fsm == 3;
  wire [1-1:0] read_rtl_bank_382;
  assign read_rtl_bank_382 = _stream_conv2d_4_source_22_source_ram_raddr;
  reg [1-1:0] _tmp_383;
  assign ram_w16_l512_id13_0_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_22_source_ram_renable && (_stream_conv2d_4_source_22_source_sel == 5))? _stream_conv2d_4_source_22_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id13_0_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_22_source_ram_renable && (_stream_conv2d_4_source_22_source_sel == 5))? 1'd1 : 0;
  localparam _tmp_384 = 1;
  wire [_tmp_384-1:0] _tmp_385;
  assign _tmp_385 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_22_source_ram_renable && (_stream_conv2d_4_source_22_source_sel == 5);
  reg [_tmp_384-1:0] __tmp_385_1;
  assign ram_w16_l512_id13_1_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_22_source_ram_renable && (_stream_conv2d_4_source_22_source_sel == 5))? _stream_conv2d_4_source_22_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id13_1_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_22_source_ram_renable && (_stream_conv2d_4_source_22_source_sel == 5))? 1'd1 : 0;
  localparam _tmp_386 = 1;
  wire [_tmp_386-1:0] _tmp_387;
  assign _tmp_387 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_22_source_ram_renable && (_stream_conv2d_4_source_22_source_sel == 5);
  reg [_tmp_386-1:0] __tmp_387_1;
  wire signed [16-1:0] read_rtl_rdata_388;
  wire read_rtl_rvalid_389;
  assign read_rtl_rdata_388 = (_tmp_383 == 0)? ram_w16_l512_id13_0_0_rdata : 
                              (_tmp_383 == 1)? ram_w16_l512_id13_1_0_rdata : 0;
  assign read_rtl_rvalid_389 = __tmp_385_1;
  assign _stream_conv2d_4_source_22_source_ram_rdata = (_stream_conv2d_4_source_22_source_sel == 5)? read_rtl_rdata_388 : 'hx;
  reg [16-1:0] __variable_wdata_1604;
  assign stream_conv2d_4_source_22_data = __variable_wdata_1604;
  reg [32-1:0] _stream_conv2d_4_source_22_source_pat_fsm_4;
  localparam _stream_conv2d_4_source_22_source_pat_fsm_4_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_22_source_pat_all_offset;
  assign _stream_conv2d_4_source_22_source_pat_all_offset = _stream_conv2d_4_source_22_source_offset_buf + _source_stream_conv2d_4_source_22_pat_cur_offset_0 + _source_stream_conv2d_4_source_22_pat_cur_offset_1 + _source_stream_conv2d_4_source_22_pat_cur_offset_2 + _source_stream_conv2d_4_source_22_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_23_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_23_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_23_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_23_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_23_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_23_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_23_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_23_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_23_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_23_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_23_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_23_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_23_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_23_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_23_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_23_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_23_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_23_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_23_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_23_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_23_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_23_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_23_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_23_pat_stride_buf_3;
  wire _set_flag_390;
  assign _set_flag_390 = conv2d_4_comp_fsm == 3;
  wire [1-1:0] read_rtl_bank_391;
  assign read_rtl_bank_391 = _stream_conv2d_4_source_23_source_ram_raddr;
  reg [1-1:0] _tmp_392;
  assign ram_w16_l512_id14_0_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_23_source_ram_renable && (_stream_conv2d_4_source_23_source_sel == 6))? _stream_conv2d_4_source_23_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id14_0_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_23_source_ram_renable && (_stream_conv2d_4_source_23_source_sel == 6))? 1'd1 : 0;
  localparam _tmp_393 = 1;
  wire [_tmp_393-1:0] _tmp_394;
  assign _tmp_394 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_23_source_ram_renable && (_stream_conv2d_4_source_23_source_sel == 6);
  reg [_tmp_393-1:0] __tmp_394_1;
  assign ram_w16_l512_id14_1_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_23_source_ram_renable && (_stream_conv2d_4_source_23_source_sel == 6))? _stream_conv2d_4_source_23_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id14_1_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_23_source_ram_renable && (_stream_conv2d_4_source_23_source_sel == 6))? 1'd1 : 0;
  localparam _tmp_395 = 1;
  wire [_tmp_395-1:0] _tmp_396;
  assign _tmp_396 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_23_source_ram_renable && (_stream_conv2d_4_source_23_source_sel == 6);
  reg [_tmp_395-1:0] __tmp_396_1;
  wire signed [16-1:0] read_rtl_rdata_397;
  wire read_rtl_rvalid_398;
  assign read_rtl_rdata_397 = (_tmp_392 == 0)? ram_w16_l512_id14_0_0_rdata : 
                              (_tmp_392 == 1)? ram_w16_l512_id14_1_0_rdata : 0;
  assign read_rtl_rvalid_398 = __tmp_394_1;
  assign _stream_conv2d_4_source_23_source_ram_rdata = (_stream_conv2d_4_source_23_source_sel == 6)? read_rtl_rdata_397 : 'hx;
  reg [16-1:0] __variable_wdata_1605;
  assign stream_conv2d_4_source_23_data = __variable_wdata_1605;
  reg [32-1:0] _stream_conv2d_4_source_23_source_pat_fsm_5;
  localparam _stream_conv2d_4_source_23_source_pat_fsm_5_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_23_source_pat_all_offset;
  assign _stream_conv2d_4_source_23_source_pat_all_offset = _stream_conv2d_4_source_23_source_offset_buf + _source_stream_conv2d_4_source_23_pat_cur_offset_0 + _source_stream_conv2d_4_source_23_pat_cur_offset_1 + _source_stream_conv2d_4_source_23_pat_cur_offset_2 + _source_stream_conv2d_4_source_23_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_24_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_24_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_24_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_24_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_24_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_24_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_24_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_24_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_24_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_24_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_24_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_24_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_24_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_24_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_24_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_24_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_24_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_24_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_24_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_24_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_24_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_24_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_24_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_24_pat_stride_buf_3;
  wire _set_flag_399;
  assign _set_flag_399 = conv2d_4_comp_fsm == 3;
  wire [1-1:0] read_rtl_bank_400;
  assign read_rtl_bank_400 = _stream_conv2d_4_source_24_source_ram_raddr;
  reg [1-1:0] _tmp_401;
  assign ram_w16_l512_id15_0_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_24_source_ram_renable && (_stream_conv2d_4_source_24_source_sel == 7))? _stream_conv2d_4_source_24_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id15_0_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_24_source_ram_renable && (_stream_conv2d_4_source_24_source_sel == 7))? 1'd1 : 0;
  localparam _tmp_402 = 1;
  wire [_tmp_402-1:0] _tmp_403;
  assign _tmp_403 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_24_source_ram_renable && (_stream_conv2d_4_source_24_source_sel == 7);
  reg [_tmp_402-1:0] __tmp_403_1;
  assign ram_w16_l512_id15_1_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_24_source_ram_renable && (_stream_conv2d_4_source_24_source_sel == 7))? _stream_conv2d_4_source_24_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id15_1_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_24_source_ram_renable && (_stream_conv2d_4_source_24_source_sel == 7))? 1'd1 : 0;
  localparam _tmp_404 = 1;
  wire [_tmp_404-1:0] _tmp_405;
  assign _tmp_405 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_24_source_ram_renable && (_stream_conv2d_4_source_24_source_sel == 7);
  reg [_tmp_404-1:0] __tmp_405_1;
  wire signed [16-1:0] read_rtl_rdata_406;
  wire read_rtl_rvalid_407;
  assign read_rtl_rdata_406 = (_tmp_401 == 0)? ram_w16_l512_id15_0_0_rdata : 
                              (_tmp_401 == 1)? ram_w16_l512_id15_1_0_rdata : 0;
  assign read_rtl_rvalid_407 = __tmp_403_1;
  assign _stream_conv2d_4_source_24_source_ram_rdata = (_stream_conv2d_4_source_24_source_sel == 7)? read_rtl_rdata_406 : 'hx;
  reg [16-1:0] __variable_wdata_1606;
  assign stream_conv2d_4_source_24_data = __variable_wdata_1606;
  reg [32-1:0] _stream_conv2d_4_source_24_source_pat_fsm_6;
  localparam _stream_conv2d_4_source_24_source_pat_fsm_6_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_24_source_pat_all_offset;
  assign _stream_conv2d_4_source_24_source_pat_all_offset = _stream_conv2d_4_source_24_source_offset_buf + _source_stream_conv2d_4_source_24_pat_cur_offset_0 + _source_stream_conv2d_4_source_24_pat_cur_offset_1 + _source_stream_conv2d_4_source_24_pat_cur_offset_2 + _source_stream_conv2d_4_source_24_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_25_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_25_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_25_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_25_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_25_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_25_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_25_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_25_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_25_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_25_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_25_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_25_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_25_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_25_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_25_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_25_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_25_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_25_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_25_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_25_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_25_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_25_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_25_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_25_pat_stride_buf_3;
  wire _set_flag_408;
  assign _set_flag_408 = conv2d_4_comp_fsm == 3;
  wire [1-1:0] read_rtl_bank_409;
  assign read_rtl_bank_409 = _stream_conv2d_4_source_25_source_ram_raddr;
  reg [1-1:0] _tmp_410;
  assign ram_w16_l512_id16_0_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_25_source_ram_renable && (_stream_conv2d_4_source_25_source_sel == 8))? _stream_conv2d_4_source_25_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id16_0_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_25_source_ram_renable && (_stream_conv2d_4_source_25_source_sel == 8))? 1'd1 : 0;
  localparam _tmp_411 = 1;
  wire [_tmp_411-1:0] _tmp_412;
  assign _tmp_412 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_25_source_ram_renable && (_stream_conv2d_4_source_25_source_sel == 8);
  reg [_tmp_411-1:0] __tmp_412_1;
  assign ram_w16_l512_id16_1_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_25_source_ram_renable && (_stream_conv2d_4_source_25_source_sel == 8))? _stream_conv2d_4_source_25_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id16_1_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_25_source_ram_renable && (_stream_conv2d_4_source_25_source_sel == 8))? 1'd1 : 0;
  localparam _tmp_413 = 1;
  wire [_tmp_413-1:0] _tmp_414;
  assign _tmp_414 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_25_source_ram_renable && (_stream_conv2d_4_source_25_source_sel == 8);
  reg [_tmp_413-1:0] __tmp_414_1;
  wire signed [16-1:0] read_rtl_rdata_415;
  wire read_rtl_rvalid_416;
  assign read_rtl_rdata_415 = (_tmp_410 == 0)? ram_w16_l512_id16_0_0_rdata : 
                              (_tmp_410 == 1)? ram_w16_l512_id16_1_0_rdata : 0;
  assign read_rtl_rvalid_416 = __tmp_412_1;
  assign _stream_conv2d_4_source_25_source_ram_rdata = (_stream_conv2d_4_source_25_source_sel == 8)? read_rtl_rdata_415 : 'hx;
  reg [16-1:0] __variable_wdata_1607;
  assign stream_conv2d_4_source_25_data = __variable_wdata_1607;
  reg [32-1:0] _stream_conv2d_4_source_25_source_pat_fsm_7;
  localparam _stream_conv2d_4_source_25_source_pat_fsm_7_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_25_source_pat_all_offset;
  assign _stream_conv2d_4_source_25_source_pat_all_offset = _stream_conv2d_4_source_25_source_offset_buf + _source_stream_conv2d_4_source_25_pat_cur_offset_0 + _source_stream_conv2d_4_source_25_pat_cur_offset_1 + _source_stream_conv2d_4_source_25_pat_cur_offset_2 + _source_stream_conv2d_4_source_25_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_26_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_26_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_26_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_26_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_26_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_26_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_26_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_26_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_26_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_26_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_26_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_26_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_26_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_26_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_26_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_26_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_26_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_26_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_26_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_26_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_26_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_26_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_26_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_26_pat_stride_buf_3;
  wire _set_flag_417;
  assign _set_flag_417 = conv2d_4_comp_fsm == 3;
  wire [1-1:0] read_rtl_bank_418;
  assign read_rtl_bank_418 = _stream_conv2d_4_source_26_source_ram_raddr;
  reg [1-1:0] _tmp_419;
  assign ram_w16_l512_id17_0_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_26_source_ram_renable && (_stream_conv2d_4_source_26_source_sel == 9))? _stream_conv2d_4_source_26_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id17_0_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_26_source_ram_renable && (_stream_conv2d_4_source_26_source_sel == 9))? 1'd1 : 0;
  localparam _tmp_420 = 1;
  wire [_tmp_420-1:0] _tmp_421;
  assign _tmp_421 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_26_source_ram_renable && (_stream_conv2d_4_source_26_source_sel == 9);
  reg [_tmp_420-1:0] __tmp_421_1;
  assign ram_w16_l512_id17_1_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_26_source_ram_renable && (_stream_conv2d_4_source_26_source_sel == 9))? _stream_conv2d_4_source_26_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id17_1_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_26_source_ram_renable && (_stream_conv2d_4_source_26_source_sel == 9))? 1'd1 : 0;
  localparam _tmp_422 = 1;
  wire [_tmp_422-1:0] _tmp_423;
  assign _tmp_423 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_26_source_ram_renable && (_stream_conv2d_4_source_26_source_sel == 9);
  reg [_tmp_422-1:0] __tmp_423_1;
  wire signed [16-1:0] read_rtl_rdata_424;
  wire read_rtl_rvalid_425;
  assign read_rtl_rdata_424 = (_tmp_419 == 0)? ram_w16_l512_id17_0_0_rdata : 
                              (_tmp_419 == 1)? ram_w16_l512_id17_1_0_rdata : 0;
  assign read_rtl_rvalid_425 = __tmp_421_1;
  assign _stream_conv2d_4_source_26_source_ram_rdata = (_stream_conv2d_4_source_26_source_sel == 9)? read_rtl_rdata_424 : 'hx;
  reg [16-1:0] __variable_wdata_1608;
  assign stream_conv2d_4_source_26_data = __variable_wdata_1608;
  reg [32-1:0] _stream_conv2d_4_source_26_source_pat_fsm_8;
  localparam _stream_conv2d_4_source_26_source_pat_fsm_8_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_26_source_pat_all_offset;
  assign _stream_conv2d_4_source_26_source_pat_all_offset = _stream_conv2d_4_source_26_source_offset_buf + _source_stream_conv2d_4_source_26_pat_cur_offset_0 + _source_stream_conv2d_4_source_26_pat_cur_offset_1 + _source_stream_conv2d_4_source_26_pat_cur_offset_2 + _source_stream_conv2d_4_source_26_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_27_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_27_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_27_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_27_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_27_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_27_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_27_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_27_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_27_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_27_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_27_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_27_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_27_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_27_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_27_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_27_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_27_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_27_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_27_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_27_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_27_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_27_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_27_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_27_pat_stride_buf_3;
  wire _set_flag_426;
  assign _set_flag_426 = conv2d_4_comp_fsm == 3;
  wire [1-1:0] read_rtl_bank_427;
  assign read_rtl_bank_427 = _stream_conv2d_4_source_27_source_ram_raddr;
  reg [1-1:0] _tmp_428;
  assign ram_w16_l512_id18_0_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_27_source_ram_renable && (_stream_conv2d_4_source_27_source_sel == 10))? _stream_conv2d_4_source_27_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id18_0_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_27_source_ram_renable && (_stream_conv2d_4_source_27_source_sel == 10))? 1'd1 : 0;
  localparam _tmp_429 = 1;
  wire [_tmp_429-1:0] _tmp_430;
  assign _tmp_430 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_27_source_ram_renable && (_stream_conv2d_4_source_27_source_sel == 10);
  reg [_tmp_429-1:0] __tmp_430_1;
  assign ram_w16_l512_id18_1_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_27_source_ram_renable && (_stream_conv2d_4_source_27_source_sel == 10))? _stream_conv2d_4_source_27_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id18_1_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_27_source_ram_renable && (_stream_conv2d_4_source_27_source_sel == 10))? 1'd1 : 0;
  localparam _tmp_431 = 1;
  wire [_tmp_431-1:0] _tmp_432;
  assign _tmp_432 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_27_source_ram_renable && (_stream_conv2d_4_source_27_source_sel == 10);
  reg [_tmp_431-1:0] __tmp_432_1;
  wire signed [16-1:0] read_rtl_rdata_433;
  wire read_rtl_rvalid_434;
  assign read_rtl_rdata_433 = (_tmp_428 == 0)? ram_w16_l512_id18_0_0_rdata : 
                              (_tmp_428 == 1)? ram_w16_l512_id18_1_0_rdata : 0;
  assign read_rtl_rvalid_434 = __tmp_430_1;
  assign _stream_conv2d_4_source_27_source_ram_rdata = (_stream_conv2d_4_source_27_source_sel == 10)? read_rtl_rdata_433 : 'hx;
  reg [16-1:0] __variable_wdata_1609;
  assign stream_conv2d_4_source_27_data = __variable_wdata_1609;
  reg [32-1:0] _stream_conv2d_4_source_27_source_pat_fsm_9;
  localparam _stream_conv2d_4_source_27_source_pat_fsm_9_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_27_source_pat_all_offset;
  assign _stream_conv2d_4_source_27_source_pat_all_offset = _stream_conv2d_4_source_27_source_offset_buf + _source_stream_conv2d_4_source_27_pat_cur_offset_0 + _source_stream_conv2d_4_source_27_pat_cur_offset_1 + _source_stream_conv2d_4_source_27_pat_cur_offset_2 + _source_stream_conv2d_4_source_27_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_28_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_28_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_28_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_28_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_28_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_28_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_28_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_28_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_28_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_28_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_28_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_28_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_28_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_28_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_28_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_28_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_28_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_28_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_28_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_28_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_28_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_28_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_28_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_28_pat_stride_buf_3;
  wire _set_flag_435;
  assign _set_flag_435 = conv2d_4_comp_fsm == 3;
  wire [1-1:0] read_rtl_bank_436;
  assign read_rtl_bank_436 = _stream_conv2d_4_source_28_source_ram_raddr;
  reg [1-1:0] _tmp_437;
  assign ram_w16_l512_id19_0_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_28_source_ram_renable && (_stream_conv2d_4_source_28_source_sel == 11))? _stream_conv2d_4_source_28_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id19_0_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_28_source_ram_renable && (_stream_conv2d_4_source_28_source_sel == 11))? 1'd1 : 0;
  localparam _tmp_438 = 1;
  wire [_tmp_438-1:0] _tmp_439;
  assign _tmp_439 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_28_source_ram_renable && (_stream_conv2d_4_source_28_source_sel == 11);
  reg [_tmp_438-1:0] __tmp_439_1;
  assign ram_w16_l512_id19_1_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_28_source_ram_renable && (_stream_conv2d_4_source_28_source_sel == 11))? _stream_conv2d_4_source_28_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id19_1_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_28_source_ram_renable && (_stream_conv2d_4_source_28_source_sel == 11))? 1'd1 : 0;
  localparam _tmp_440 = 1;
  wire [_tmp_440-1:0] _tmp_441;
  assign _tmp_441 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_28_source_ram_renable && (_stream_conv2d_4_source_28_source_sel == 11);
  reg [_tmp_440-1:0] __tmp_441_1;
  wire signed [16-1:0] read_rtl_rdata_442;
  wire read_rtl_rvalid_443;
  assign read_rtl_rdata_442 = (_tmp_437 == 0)? ram_w16_l512_id19_0_0_rdata : 
                              (_tmp_437 == 1)? ram_w16_l512_id19_1_0_rdata : 0;
  assign read_rtl_rvalid_443 = __tmp_439_1;
  assign _stream_conv2d_4_source_28_source_ram_rdata = (_stream_conv2d_4_source_28_source_sel == 11)? read_rtl_rdata_442 : 'hx;
  reg [16-1:0] __variable_wdata_1610;
  assign stream_conv2d_4_source_28_data = __variable_wdata_1610;
  reg [32-1:0] _stream_conv2d_4_source_28_source_pat_fsm_10;
  localparam _stream_conv2d_4_source_28_source_pat_fsm_10_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_28_source_pat_all_offset;
  assign _stream_conv2d_4_source_28_source_pat_all_offset = _stream_conv2d_4_source_28_source_offset_buf + _source_stream_conv2d_4_source_28_pat_cur_offset_0 + _source_stream_conv2d_4_source_28_pat_cur_offset_1 + _source_stream_conv2d_4_source_28_pat_cur_offset_2 + _source_stream_conv2d_4_source_28_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_29_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_29_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_29_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_29_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_29_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_29_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_29_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_29_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_29_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_29_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_29_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_29_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_29_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_29_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_29_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_29_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_29_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_29_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_29_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_29_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_29_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_29_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_29_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_29_pat_stride_buf_3;
  wire _set_flag_444;
  assign _set_flag_444 = conv2d_4_comp_fsm == 3;
  wire [1-1:0] read_rtl_bank_445;
  assign read_rtl_bank_445 = _stream_conv2d_4_source_29_source_ram_raddr;
  reg [1-1:0] _tmp_446;
  localparam _tmp_447 = 1;
  wire [_tmp_447-1:0] _tmp_448;
  assign _tmp_448 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_29_source_ram_renable && (_stream_conv2d_4_source_29_source_sel == 12);
  reg [_tmp_447-1:0] __tmp_448_1;
  localparam _tmp_449 = 1;
  wire [_tmp_449-1:0] _tmp_450;
  assign _tmp_450 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_29_source_ram_renable && (_stream_conv2d_4_source_29_source_sel == 12);
  reg [_tmp_449-1:0] __tmp_450_1;
  wire signed [16-1:0] read_rtl_rdata_451;
  wire read_rtl_rvalid_452;
  assign read_rtl_rdata_451 = (_tmp_446 == 0)? ram_w16_l512_id0_0_0_rdata : 
                              (_tmp_446 == 1)? ram_w16_l512_id0_1_0_rdata : 0;
  assign read_rtl_rvalid_452 = __tmp_448_1;
  assign _stream_conv2d_4_source_29_source_ram_rdata = (_stream_conv2d_4_source_29_source_sel == 12)? read_rtl_rdata_451 : 'hx;
  reg [16-1:0] __variable_wdata_1836;
  assign stream_conv2d_4_source_29_data = __variable_wdata_1836;
  reg [32-1:0] _stream_conv2d_4_source_29_source_pat_fsm_11;
  localparam _stream_conv2d_4_source_29_source_pat_fsm_11_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_29_source_pat_all_offset;
  assign _stream_conv2d_4_source_29_source_pat_all_offset = _stream_conv2d_4_source_29_source_offset_buf + _source_stream_conv2d_4_source_29_pat_cur_offset_0 + _source_stream_conv2d_4_source_29_pat_cur_offset_1 + _source_stream_conv2d_4_source_29_pat_cur_offset_2 + _source_stream_conv2d_4_source_29_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_30_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_30_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_30_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_30_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_30_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_30_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_30_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_30_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_30_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_30_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_30_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_30_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_30_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_30_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_30_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_30_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_30_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_30_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_30_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_30_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_30_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_30_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_30_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_30_pat_stride_buf_3;
  wire _set_flag_453;
  assign _set_flag_453 = conv2d_4_comp_fsm == 3;
  wire [1-1:0] read_rtl_bank_454;
  assign read_rtl_bank_454 = _stream_conv2d_4_source_30_source_ram_raddr;
  reg [1-1:0] _tmp_455;
  localparam _tmp_456 = 1;
  wire [_tmp_456-1:0] _tmp_457;
  assign _tmp_457 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_30_source_ram_renable && (_stream_conv2d_4_source_30_source_sel == 13);
  reg [_tmp_456-1:0] __tmp_457_1;
  localparam _tmp_458 = 1;
  wire [_tmp_458-1:0] _tmp_459;
  assign _tmp_459 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_30_source_ram_renable && (_stream_conv2d_4_source_30_source_sel == 13);
  reg [_tmp_458-1:0] __tmp_459_1;
  wire signed [16-1:0] read_rtl_rdata_460;
  wire read_rtl_rvalid_461;
  assign read_rtl_rdata_460 = (_tmp_455 == 0)? ram_w16_l512_id1_0_0_rdata : 
                              (_tmp_455 == 1)? ram_w16_l512_id1_1_0_rdata : 0;
  assign read_rtl_rvalid_461 = __tmp_457_1;
  assign _stream_conv2d_4_source_30_source_ram_rdata = (_stream_conv2d_4_source_30_source_sel == 13)? read_rtl_rdata_460 : 'hx;
  reg [16-1:0] __variable_wdata_1837;
  assign stream_conv2d_4_source_30_data = __variable_wdata_1837;
  reg [32-1:0] _stream_conv2d_4_source_30_source_pat_fsm_12;
  localparam _stream_conv2d_4_source_30_source_pat_fsm_12_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_30_source_pat_all_offset;
  assign _stream_conv2d_4_source_30_source_pat_all_offset = _stream_conv2d_4_source_30_source_offset_buf + _source_stream_conv2d_4_source_30_pat_cur_offset_0 + _source_stream_conv2d_4_source_30_pat_cur_offset_1 + _source_stream_conv2d_4_source_30_pat_cur_offset_2 + _source_stream_conv2d_4_source_30_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_31_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_31_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_31_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_31_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_31_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_31_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_31_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_31_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_31_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_31_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_31_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_31_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_31_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_31_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_31_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_31_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_31_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_31_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_31_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_31_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_31_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_31_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_31_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_31_pat_stride_buf_3;
  wire _set_flag_462;
  assign _set_flag_462 = conv2d_4_comp_fsm == 3;
  wire [1-1:0] read_rtl_bank_463;
  assign read_rtl_bank_463 = _stream_conv2d_4_source_31_source_ram_raddr;
  reg [1-1:0] _tmp_464;
  localparam _tmp_465 = 1;
  wire [_tmp_465-1:0] _tmp_466;
  assign _tmp_466 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_31_source_ram_renable && (_stream_conv2d_4_source_31_source_sel == 14);
  reg [_tmp_465-1:0] __tmp_466_1;
  localparam _tmp_467 = 1;
  wire [_tmp_467-1:0] _tmp_468;
  assign _tmp_468 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_31_source_ram_renable && (_stream_conv2d_4_source_31_source_sel == 14);
  reg [_tmp_467-1:0] __tmp_468_1;
  wire signed [16-1:0] read_rtl_rdata_469;
  wire read_rtl_rvalid_470;
  assign read_rtl_rdata_469 = (_tmp_464 == 0)? ram_w16_l512_id2_0_0_rdata : 
                              (_tmp_464 == 1)? ram_w16_l512_id2_1_0_rdata : 0;
  assign read_rtl_rvalid_470 = __tmp_466_1;
  assign _stream_conv2d_4_source_31_source_ram_rdata = (_stream_conv2d_4_source_31_source_sel == 14)? read_rtl_rdata_469 : 'hx;
  reg [16-1:0] __variable_wdata_1838;
  assign stream_conv2d_4_source_31_data = __variable_wdata_1838;
  reg [32-1:0] _stream_conv2d_4_source_31_source_pat_fsm_13;
  localparam _stream_conv2d_4_source_31_source_pat_fsm_13_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_31_source_pat_all_offset;
  assign _stream_conv2d_4_source_31_source_pat_all_offset = _stream_conv2d_4_source_31_source_offset_buf + _source_stream_conv2d_4_source_31_pat_cur_offset_0 + _source_stream_conv2d_4_source_31_pat_cur_offset_1 + _source_stream_conv2d_4_source_31_pat_cur_offset_2 + _source_stream_conv2d_4_source_31_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_32_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_32_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_32_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_32_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_32_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_32_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_32_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_32_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_32_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_32_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_32_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_32_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_32_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_32_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_32_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_32_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_32_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_32_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_32_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_32_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_32_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_32_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_32_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_32_pat_stride_buf_3;
  wire _set_flag_471;
  assign _set_flag_471 = conv2d_4_comp_fsm == 3;
  wire [1-1:0] read_rtl_bank_472;
  assign read_rtl_bank_472 = _stream_conv2d_4_source_32_source_ram_raddr;
  reg [1-1:0] _tmp_473;
  assign ram_w16_l512_id3_0_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_32_source_ram_renable && (_stream_conv2d_4_source_32_source_sel == 15))? _stream_conv2d_4_source_32_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id3_0_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_32_source_ram_renable && (_stream_conv2d_4_source_32_source_sel == 15))? 1'd1 : 0;
  localparam _tmp_474 = 1;
  wire [_tmp_474-1:0] _tmp_475;
  assign _tmp_475 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_32_source_ram_renable && (_stream_conv2d_4_source_32_source_sel == 15);
  reg [_tmp_474-1:0] __tmp_475_1;
  assign ram_w16_l512_id3_1_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_32_source_ram_renable && (_stream_conv2d_4_source_32_source_sel == 15))? _stream_conv2d_4_source_32_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id3_1_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_32_source_ram_renable && (_stream_conv2d_4_source_32_source_sel == 15))? 1'd1 : 0;
  localparam _tmp_476 = 1;
  wire [_tmp_476-1:0] _tmp_477;
  assign _tmp_477 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_32_source_ram_renable && (_stream_conv2d_4_source_32_source_sel == 15);
  reg [_tmp_476-1:0] __tmp_477_1;
  wire signed [16-1:0] read_rtl_rdata_478;
  wire read_rtl_rvalid_479;
  assign read_rtl_rdata_478 = (_tmp_473 == 0)? ram_w16_l512_id3_0_0_rdata : 
                              (_tmp_473 == 1)? ram_w16_l512_id3_1_0_rdata : 0;
  assign read_rtl_rvalid_479 = __tmp_475_1;
  assign _stream_conv2d_4_source_32_source_ram_rdata = (_stream_conv2d_4_source_32_source_sel == 15)? read_rtl_rdata_478 : 'hx;
  reg [16-1:0] __variable_wdata_1839;
  assign stream_conv2d_4_source_32_data = __variable_wdata_1839;
  reg [32-1:0] _stream_conv2d_4_source_32_source_pat_fsm_14;
  localparam _stream_conv2d_4_source_32_source_pat_fsm_14_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_32_source_pat_all_offset;
  assign _stream_conv2d_4_source_32_source_pat_all_offset = _stream_conv2d_4_source_32_source_offset_buf + _source_stream_conv2d_4_source_32_pat_cur_offset_0 + _source_stream_conv2d_4_source_32_pat_cur_offset_1 + _source_stream_conv2d_4_source_32_pat_cur_offset_2 + _source_stream_conv2d_4_source_32_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_33_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_33_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_33_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_33_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_33_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_33_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_33_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_33_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_33_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_33_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_33_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_33_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_33_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_33_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_33_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_33_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_33_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_33_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_33_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_33_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_33_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_33_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_33_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_33_pat_stride_buf_3;
  wire _set_flag_480;
  assign _set_flag_480 = conv2d_4_comp_fsm == 3;
  wire [1-1:0] read_rtl_bank_481;
  assign read_rtl_bank_481 = _stream_conv2d_4_source_33_source_ram_raddr;
  reg [1-1:0] _tmp_482;
  assign ram_w16_l512_id4_0_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_33_source_ram_renable && (_stream_conv2d_4_source_33_source_sel == 16))? _stream_conv2d_4_source_33_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id4_0_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_33_source_ram_renable && (_stream_conv2d_4_source_33_source_sel == 16))? 1'd1 : 0;
  localparam _tmp_483 = 1;
  wire [_tmp_483-1:0] _tmp_484;
  assign _tmp_484 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_33_source_ram_renable && (_stream_conv2d_4_source_33_source_sel == 16);
  reg [_tmp_483-1:0] __tmp_484_1;
  assign ram_w16_l512_id4_1_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_33_source_ram_renable && (_stream_conv2d_4_source_33_source_sel == 16))? _stream_conv2d_4_source_33_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id4_1_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_33_source_ram_renable && (_stream_conv2d_4_source_33_source_sel == 16))? 1'd1 : 0;
  localparam _tmp_485 = 1;
  wire [_tmp_485-1:0] _tmp_486;
  assign _tmp_486 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_33_source_ram_renable && (_stream_conv2d_4_source_33_source_sel == 16);
  reg [_tmp_485-1:0] __tmp_486_1;
  wire signed [16-1:0] read_rtl_rdata_487;
  wire read_rtl_rvalid_488;
  assign read_rtl_rdata_487 = (_tmp_482 == 0)? ram_w16_l512_id4_0_0_rdata : 
                              (_tmp_482 == 1)? ram_w16_l512_id4_1_0_rdata : 0;
  assign read_rtl_rvalid_488 = __tmp_484_1;
  assign _stream_conv2d_4_source_33_source_ram_rdata = (_stream_conv2d_4_source_33_source_sel == 16)? read_rtl_rdata_487 : 'hx;
  reg [16-1:0] __variable_wdata_1840;
  assign stream_conv2d_4_source_33_data = __variable_wdata_1840;
  reg [32-1:0] _stream_conv2d_4_source_33_source_pat_fsm_15;
  localparam _stream_conv2d_4_source_33_source_pat_fsm_15_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_33_source_pat_all_offset;
  assign _stream_conv2d_4_source_33_source_pat_all_offset = _stream_conv2d_4_source_33_source_offset_buf + _source_stream_conv2d_4_source_33_pat_cur_offset_0 + _source_stream_conv2d_4_source_33_pat_cur_offset_1 + _source_stream_conv2d_4_source_33_pat_cur_offset_2 + _source_stream_conv2d_4_source_33_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_34_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_34_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_34_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_34_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_34_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_34_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_34_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_34_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_34_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_34_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_34_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_34_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_34_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_34_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_34_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_34_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_34_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_34_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_34_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_34_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_34_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_34_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_34_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_34_pat_stride_buf_3;
  wire _set_flag_489;
  assign _set_flag_489 = conv2d_4_comp_fsm == 3;
  wire [1-1:0] read_rtl_bank_490;
  assign read_rtl_bank_490 = _stream_conv2d_4_source_34_source_ram_raddr;
  reg [1-1:0] _tmp_491;
  assign ram_w16_l512_id5_0_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_34_source_ram_renable && (_stream_conv2d_4_source_34_source_sel == 17))? _stream_conv2d_4_source_34_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id5_0_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_34_source_ram_renable && (_stream_conv2d_4_source_34_source_sel == 17))? 1'd1 : 0;
  localparam _tmp_492 = 1;
  wire [_tmp_492-1:0] _tmp_493;
  assign _tmp_493 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_34_source_ram_renable && (_stream_conv2d_4_source_34_source_sel == 17);
  reg [_tmp_492-1:0] __tmp_493_1;
  assign ram_w16_l512_id5_1_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_34_source_ram_renable && (_stream_conv2d_4_source_34_source_sel == 17))? _stream_conv2d_4_source_34_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id5_1_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_34_source_ram_renable && (_stream_conv2d_4_source_34_source_sel == 17))? 1'd1 : 0;
  localparam _tmp_494 = 1;
  wire [_tmp_494-1:0] _tmp_495;
  assign _tmp_495 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_34_source_ram_renable && (_stream_conv2d_4_source_34_source_sel == 17);
  reg [_tmp_494-1:0] __tmp_495_1;
  wire signed [16-1:0] read_rtl_rdata_496;
  wire read_rtl_rvalid_497;
  assign read_rtl_rdata_496 = (_tmp_491 == 0)? ram_w16_l512_id5_0_0_rdata : 
                              (_tmp_491 == 1)? ram_w16_l512_id5_1_0_rdata : 0;
  assign read_rtl_rvalid_497 = __tmp_493_1;
  assign _stream_conv2d_4_source_34_source_ram_rdata = (_stream_conv2d_4_source_34_source_sel == 17)? read_rtl_rdata_496 : 'hx;
  reg [16-1:0] __variable_wdata_1841;
  assign stream_conv2d_4_source_34_data = __variable_wdata_1841;
  reg [32-1:0] _stream_conv2d_4_source_34_source_pat_fsm_16;
  localparam _stream_conv2d_4_source_34_source_pat_fsm_16_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_34_source_pat_all_offset;
  assign _stream_conv2d_4_source_34_source_pat_all_offset = _stream_conv2d_4_source_34_source_offset_buf + _source_stream_conv2d_4_source_34_pat_cur_offset_0 + _source_stream_conv2d_4_source_34_pat_cur_offset_1 + _source_stream_conv2d_4_source_34_pat_cur_offset_2 + _source_stream_conv2d_4_source_34_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_35_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_35_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_35_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_35_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_35_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_35_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_35_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_35_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_35_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_35_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_35_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_35_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_35_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_35_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_35_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_35_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_35_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_35_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_35_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_35_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_35_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_35_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_35_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_35_pat_stride_buf_3;
  wire _set_flag_498;
  assign _set_flag_498 = conv2d_4_comp_fsm == 3;
  wire [1-1:0] read_rtl_bank_499;
  assign read_rtl_bank_499 = _stream_conv2d_4_source_35_source_ram_raddr;
  reg [1-1:0] _tmp_500;
  assign ram_w16_l512_id6_0_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_35_source_ram_renable && (_stream_conv2d_4_source_35_source_sel == 18))? _stream_conv2d_4_source_35_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id6_0_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_35_source_ram_renable && (_stream_conv2d_4_source_35_source_sel == 18))? 1'd1 : 0;
  localparam _tmp_501 = 1;
  wire [_tmp_501-1:0] _tmp_502;
  assign _tmp_502 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_35_source_ram_renable && (_stream_conv2d_4_source_35_source_sel == 18);
  reg [_tmp_501-1:0] __tmp_502_1;
  assign ram_w16_l512_id6_1_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_35_source_ram_renable && (_stream_conv2d_4_source_35_source_sel == 18))? _stream_conv2d_4_source_35_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id6_1_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_35_source_ram_renable && (_stream_conv2d_4_source_35_source_sel == 18))? 1'd1 : 0;
  localparam _tmp_503 = 1;
  wire [_tmp_503-1:0] _tmp_504;
  assign _tmp_504 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_35_source_ram_renable && (_stream_conv2d_4_source_35_source_sel == 18);
  reg [_tmp_503-1:0] __tmp_504_1;
  wire signed [16-1:0] read_rtl_rdata_505;
  wire read_rtl_rvalid_506;
  assign read_rtl_rdata_505 = (_tmp_500 == 0)? ram_w16_l512_id6_0_0_rdata : 
                              (_tmp_500 == 1)? ram_w16_l512_id6_1_0_rdata : 0;
  assign read_rtl_rvalid_506 = __tmp_502_1;
  assign _stream_conv2d_4_source_35_source_ram_rdata = (_stream_conv2d_4_source_35_source_sel == 18)? read_rtl_rdata_505 : 'hx;
  reg [16-1:0] __variable_wdata_1842;
  assign stream_conv2d_4_source_35_data = __variable_wdata_1842;
  reg [32-1:0] _stream_conv2d_4_source_35_source_pat_fsm_17;
  localparam _stream_conv2d_4_source_35_source_pat_fsm_17_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_35_source_pat_all_offset;
  assign _stream_conv2d_4_source_35_source_pat_all_offset = _stream_conv2d_4_source_35_source_offset_buf + _source_stream_conv2d_4_source_35_pat_cur_offset_0 + _source_stream_conv2d_4_source_35_pat_cur_offset_1 + _source_stream_conv2d_4_source_35_pat_cur_offset_2 + _source_stream_conv2d_4_source_35_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_36_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_36_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_36_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_36_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_36_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_36_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_36_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_36_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_36_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_36_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_36_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_36_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_36_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_36_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_36_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_36_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_36_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_36_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_36_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_36_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_36_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_36_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_36_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_36_pat_stride_buf_3;
  wire _set_flag_507;
  assign _set_flag_507 = conv2d_4_comp_fsm == 3;
  wire [1-1:0] read_rtl_bank_508;
  assign read_rtl_bank_508 = _stream_conv2d_4_source_36_source_ram_raddr;
  reg [1-1:0] _tmp_509;
  assign ram_w16_l512_id7_0_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_36_source_ram_renable && (_stream_conv2d_4_source_36_source_sel == 19))? _stream_conv2d_4_source_36_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id7_0_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_36_source_ram_renable && (_stream_conv2d_4_source_36_source_sel == 19))? 1'd1 : 0;
  localparam _tmp_510 = 1;
  wire [_tmp_510-1:0] _tmp_511;
  assign _tmp_511 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_36_source_ram_renable && (_stream_conv2d_4_source_36_source_sel == 19);
  reg [_tmp_510-1:0] __tmp_511_1;
  assign ram_w16_l512_id7_1_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_36_source_ram_renable && (_stream_conv2d_4_source_36_source_sel == 19))? _stream_conv2d_4_source_36_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id7_1_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_36_source_ram_renable && (_stream_conv2d_4_source_36_source_sel == 19))? 1'd1 : 0;
  localparam _tmp_512 = 1;
  wire [_tmp_512-1:0] _tmp_513;
  assign _tmp_513 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_36_source_ram_renable && (_stream_conv2d_4_source_36_source_sel == 19);
  reg [_tmp_512-1:0] __tmp_513_1;
  wire signed [16-1:0] read_rtl_rdata_514;
  wire read_rtl_rvalid_515;
  assign read_rtl_rdata_514 = (_tmp_509 == 0)? ram_w16_l512_id7_0_0_rdata : 
                              (_tmp_509 == 1)? ram_w16_l512_id7_1_0_rdata : 0;
  assign read_rtl_rvalid_515 = __tmp_511_1;
  assign _stream_conv2d_4_source_36_source_ram_rdata = (_stream_conv2d_4_source_36_source_sel == 19)? read_rtl_rdata_514 : 'hx;
  reg [16-1:0] __variable_wdata_1843;
  assign stream_conv2d_4_source_36_data = __variable_wdata_1843;
  reg [32-1:0] _stream_conv2d_4_source_36_source_pat_fsm_18;
  localparam _stream_conv2d_4_source_36_source_pat_fsm_18_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_36_source_pat_all_offset;
  assign _stream_conv2d_4_source_36_source_pat_all_offset = _stream_conv2d_4_source_36_source_offset_buf + _source_stream_conv2d_4_source_36_pat_cur_offset_0 + _source_stream_conv2d_4_source_36_pat_cur_offset_1 + _source_stream_conv2d_4_source_36_pat_cur_offset_2 + _source_stream_conv2d_4_source_36_pat_cur_offset_3;
  reg [32-1:0] _source_stream_conv2d_4_source_37_pat_cur_offset_0;
  reg [32-1:0] _source_stream_conv2d_4_source_37_pat_cur_offset_1;
  reg [32-1:0] _source_stream_conv2d_4_source_37_pat_cur_offset_2;
  reg [32-1:0] _source_stream_conv2d_4_source_37_pat_cur_offset_3;
  reg [33-1:0] _source_stream_conv2d_4_source_37_pat_size_0;
  reg [33-1:0] _source_stream_conv2d_4_source_37_pat_size_1;
  reg [33-1:0] _source_stream_conv2d_4_source_37_pat_size_2;
  reg [33-1:0] _source_stream_conv2d_4_source_37_pat_size_3;
  reg [32-1:0] _source_stream_conv2d_4_source_37_pat_stride_0;
  reg [32-1:0] _source_stream_conv2d_4_source_37_pat_stride_1;
  reg [32-1:0] _source_stream_conv2d_4_source_37_pat_stride_2;
  reg [32-1:0] _source_stream_conv2d_4_source_37_pat_stride_3;
  reg [33-1:0] _source_stream_conv2d_4_source_37_pat_count_0;
  reg [33-1:0] _source_stream_conv2d_4_source_37_pat_count_1;
  reg [33-1:0] _source_stream_conv2d_4_source_37_pat_count_2;
  reg [33-1:0] _source_stream_conv2d_4_source_37_pat_count_3;
  reg [33-1:0] _source_stream_conv2d_4_source_37_pat_size_buf_0;
  reg [33-1:0] _source_stream_conv2d_4_source_37_pat_size_buf_1;
  reg [33-1:0] _source_stream_conv2d_4_source_37_pat_size_buf_2;
  reg [33-1:0] _source_stream_conv2d_4_source_37_pat_size_buf_3;
  reg [32-1:0] _source_stream_conv2d_4_source_37_pat_stride_buf_0;
  reg [32-1:0] _source_stream_conv2d_4_source_37_pat_stride_buf_1;
  reg [32-1:0] _source_stream_conv2d_4_source_37_pat_stride_buf_2;
  reg [32-1:0] _source_stream_conv2d_4_source_37_pat_stride_buf_3;
  wire _set_flag_516;
  assign _set_flag_516 = conv2d_4_comp_fsm == 3;
  wire [1-1:0] read_rtl_bank_517;
  assign read_rtl_bank_517 = _stream_conv2d_4_source_37_source_ram_raddr;
  reg [1-1:0] _tmp_518;
  assign ram_w16_l512_id8_0_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_37_source_ram_renable && (_stream_conv2d_4_source_37_source_sel == 20))? _stream_conv2d_4_source_37_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id8_0_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_37_source_ram_renable && (_stream_conv2d_4_source_37_source_sel == 20))? 1'd1 : 0;
  localparam _tmp_519 = 1;
  wire [_tmp_519-1:0] _tmp_520;
  assign _tmp_520 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_37_source_ram_renable && (_stream_conv2d_4_source_37_source_sel == 20);
  reg [_tmp_519-1:0] __tmp_520_1;
  assign ram_w16_l512_id8_1_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_37_source_ram_renable && (_stream_conv2d_4_source_37_source_sel == 20))? _stream_conv2d_4_source_37_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id8_1_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_37_source_ram_renable && (_stream_conv2d_4_source_37_source_sel == 20))? 1'd1 : 0;
  localparam _tmp_521 = 1;
  wire [_tmp_521-1:0] _tmp_522;
  assign _tmp_522 = _stream_conv2d_4_stream_oready && _stream_conv2d_4_source_37_source_ram_renable && (_stream_conv2d_4_source_37_source_sel == 20);
  reg [_tmp_521-1:0] __tmp_522_1;
  wire signed [16-1:0] read_rtl_rdata_523;
  wire read_rtl_rvalid_524;
  assign read_rtl_rdata_523 = (_tmp_518 == 0)? ram_w16_l512_id8_0_0_rdata : 
                              (_tmp_518 == 1)? ram_w16_l512_id8_1_0_rdata : 0;
  assign read_rtl_rvalid_524 = __tmp_520_1;
  assign _stream_conv2d_4_source_37_source_ram_rdata = (_stream_conv2d_4_source_37_source_sel == 20)? read_rtl_rdata_523 : 'hx;
  reg [16-1:0] __variable_wdata_1844;
  assign stream_conv2d_4_source_37_data = __variable_wdata_1844;
  reg [32-1:0] _stream_conv2d_4_source_37_source_pat_fsm_19;
  localparam _stream_conv2d_4_source_37_source_pat_fsm_19_init = 0;
  wire [32-1:0] _stream_conv2d_4_source_37_source_pat_all_offset;
  assign _stream_conv2d_4_source_37_source_pat_all_offset = _stream_conv2d_4_source_37_source_offset_buf + _source_stream_conv2d_4_source_37_pat_cur_offset_0 + _source_stream_conv2d_4_source_37_pat_cur_offset_1 + _source_stream_conv2d_4_source_37_pat_cur_offset_2 + _source_stream_conv2d_4_source_37_pat_cur_offset_3;
  wire _set_flag_525;
  assign _set_flag_525 = conv2d_4_comp_fsm == 3;
  reg _tmp_526;
  reg _tmp_527;
  reg _tmp_528;
  reg _tmp_529;
  reg _tmp_530;
  reg _tmp_531;
  reg _tmp_532;
  reg _tmp_533;
  reg _tmp_534;
  reg _tmp_535;
  reg _tmp_536;
  reg _tmp_537;
  reg _tmp_538;
  reg _tmp_539;
  reg _tmp_540;
  reg _tmp_541;
  reg _tmp_542;
  reg _tmp_543;
  reg _tmp_544;
  reg _tmp_545;
  reg _tmp_546;
  reg _tmp_547;
  reg _tmp_548;
  reg _tmp_549;
  reg _tmp_550;
  reg _tmp_551;
  reg _tmp_552;
  reg _tmp_553;
  reg _tmp_554;
  reg _tmp_555;
  reg _tmp_556;
  reg _tmp_557;
  reg _tmp_558;
  localparam _tmp_559 = 33;
  wire [_tmp_559-1:0] _tmp_560;
  assign _tmp_560 = conv2d_4_stream_out_local + conv2d_4_out_page_comp_offset_buf;
  reg [_tmp_559-1:0] _tmp_561;
  reg [_tmp_559-1:0] _tmp_562;
  reg [_tmp_559-1:0] _tmp_563;
  reg [_tmp_559-1:0] _tmp_564;
  reg [_tmp_559-1:0] _tmp_565;
  reg [_tmp_559-1:0] _tmp_566;
  reg [_tmp_559-1:0] _tmp_567;
  reg [_tmp_559-1:0] _tmp_568;
  reg [_tmp_559-1:0] _tmp_569;
  reg [_tmp_559-1:0] _tmp_570;
  reg [_tmp_559-1:0] _tmp_571;
  reg [_tmp_559-1:0] _tmp_572;
  reg [_tmp_559-1:0] _tmp_573;
  reg [_tmp_559-1:0] _tmp_574;
  reg [_tmp_559-1:0] _tmp_575;
  reg [_tmp_559-1:0] _tmp_576;
  reg [_tmp_559-1:0] _tmp_577;
  reg [_tmp_559-1:0] _tmp_578;
  reg [_tmp_559-1:0] _tmp_579;
  reg [_tmp_559-1:0] _tmp_580;
  reg [_tmp_559-1:0] _tmp_581;
  reg [_tmp_559-1:0] _tmp_582;
  reg [_tmp_559-1:0] _tmp_583;
  reg [_tmp_559-1:0] _tmp_584;
  reg [_tmp_559-1:0] _tmp_585;
  reg [_tmp_559-1:0] _tmp_586;
  reg [_tmp_559-1:0] _tmp_587;
  reg [_tmp_559-1:0] _tmp_588;
  reg [_tmp_559-1:0] _tmp_589;
  reg [_tmp_559-1:0] _tmp_590;
  reg [_tmp_559-1:0] _tmp_591;
  reg [_tmp_559-1:0] _tmp_592;
  reg [_tmp_559-1:0] _tmp_593;
  reg [32-1:0] _tmp_594;
  reg [32-1:0] _tmp_595;
  reg [32-1:0] _tmp_596;
  reg [32-1:0] _tmp_597;
  reg [32-1:0] _tmp_598;
  reg [32-1:0] _tmp_599;
  reg [32-1:0] _tmp_600;
  reg [32-1:0] _tmp_601;
  reg [32-1:0] _tmp_602;
  reg [32-1:0] _tmp_603;
  reg [32-1:0] _tmp_604;
  reg [32-1:0] _tmp_605;
  reg [32-1:0] _tmp_606;
  reg [32-1:0] _tmp_607;
  reg [32-1:0] _tmp_608;
  reg [32-1:0] _tmp_609;
  reg [32-1:0] _tmp_610;
  reg [32-1:0] _tmp_611;
  reg [32-1:0] _tmp_612;
  reg [32-1:0] _tmp_613;
  reg [32-1:0] _tmp_614;
  reg [32-1:0] _tmp_615;
  reg [32-1:0] _tmp_616;
  reg [32-1:0] _tmp_617;
  reg [32-1:0] _tmp_618;
  reg [32-1:0] _tmp_619;
  reg [32-1:0] _tmp_620;
  reg [32-1:0] _tmp_621;
  reg [32-1:0] _tmp_622;
  reg [32-1:0] _tmp_623;
  reg [32-1:0] _tmp_624;
  reg [32-1:0] _tmp_625;
  reg [32-1:0] _tmp_626;
  wire [1-1:0] write_rtl_bank_627;
  assign write_rtl_bank_627 = _stream_conv2d_4_sink_50_sink_waddr;
  assign ram_w16_l512_id20_0_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_sink_50_sink_wenable && (_stream_conv2d_4_sink_50_sink_sel == 21) && (write_rtl_bank_627 == 0))? _stream_conv2d_4_sink_50_sink_waddr >> 1 : 'hx;
  assign ram_w16_l512_id20_0_0_wdata = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_sink_50_sink_wenable && (_stream_conv2d_4_sink_50_sink_sel == 21) && (write_rtl_bank_627 == 0))? _stream_conv2d_4_sink_50_sink_wdata : 'hx;
  assign ram_w16_l512_id20_0_0_wenable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_sink_50_sink_wenable && (_stream_conv2d_4_sink_50_sink_sel == 21) && (write_rtl_bank_627 == 0))? 1'd1 : 0;
  assign ram_w16_l512_id20_0_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_sink_50_sink_wenable && (_stream_conv2d_4_sink_50_sink_sel == 21) && (write_rtl_bank_627 == 0))? 1'd1 : 0;
  assign ram_w16_l512_id20_1_0_addr = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_sink_50_sink_wenable && (_stream_conv2d_4_sink_50_sink_sel == 21) && (write_rtl_bank_627 == 1))? _stream_conv2d_4_sink_50_sink_waddr >> 1 : 'hx;
  assign ram_w16_l512_id20_1_0_wdata = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_sink_50_sink_wenable && (_stream_conv2d_4_sink_50_sink_sel == 21) && (write_rtl_bank_627 == 1))? _stream_conv2d_4_sink_50_sink_wdata : 'hx;
  assign ram_w16_l512_id20_1_0_wenable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_sink_50_sink_wenable && (_stream_conv2d_4_sink_50_sink_sel == 21) && (write_rtl_bank_627 == 1))? 1'd1 : 0;
  assign ram_w16_l512_id20_1_0_enable = (_stream_conv2d_4_stream_oready && _stream_conv2d_4_sink_50_sink_wenable && (_stream_conv2d_4_sink_50_sink_sel == 21) && (write_rtl_bank_627 == 1))? 1'd1 : 0;
  reg [32-1:0] _stream_conv2d_4_sink_50_sink_fsm_20;
  localparam _stream_conv2d_4_sink_50_sink_fsm_20_init = 0;
  wire _set_flag_628;
  assign _set_flag_628 = conv2d_4_comp_fsm == 4;
  assign _stream_conv2d_4_run_flag = (_set_flag_628)? 1 : 0;
  reg _tmp_629;
  reg _tmp_630;
  reg _tmp_631;
  assign _mul_18_source_stop = _mul_18_stream_oready && 1'd0;
  reg _tmp_632;
  reg _tmp_633;
  reg _tmp_634;
  reg _tmp_635;
  reg _tmp_636;
  reg _tmp_637;
  reg _tmp_638;
  reg _tmp_639;
  reg _tmp_640;
  reg _tmp_641;
  assign _mul_18_sink_start = _tmp_641;
  reg _tmp_642;
  reg _tmp_643;
  reg _tmp_644;
  reg _tmp_645;
  reg _tmp_646;
  reg _tmp_647;
  reg _tmp_648;
  reg _tmp_649;
  reg _tmp_650;
  reg _tmp_651;
  assign _mul_18_sink_stop = _tmp_651;
  reg _tmp_652;
  reg _tmp_653;
  reg _tmp_654;
  reg _tmp_655;
  reg _tmp_656;
  reg _tmp_657;
  reg _tmp_658;
  reg _tmp_659;
  reg _tmp_660;
  reg _tmp_661;
  assign _mul_18_sink_busy = _tmp_661;
  reg _tmp_662;
  assign _mul_18_busy = _mul_18_source_busy || _mul_18_sink_busy || _mul_18_busy_reg;
  reg _tmp_663;
  reg _tmp_664;
  reg _tmp_665;
  assign _mul_19_source_stop = _mul_19_stream_oready && 1'd0;
  reg _tmp_666;
  reg _tmp_667;
  reg _tmp_668;
  reg _tmp_669;
  reg _tmp_670;
  reg _tmp_671;
  reg _tmp_672;
  reg _tmp_673;
  reg _tmp_674;
  reg _tmp_675;
  assign _mul_19_sink_start = _tmp_675;
  reg _tmp_676;
  reg _tmp_677;
  reg _tmp_678;
  reg _tmp_679;
  reg _tmp_680;
  reg _tmp_681;
  reg _tmp_682;
  reg _tmp_683;
  reg _tmp_684;
  reg _tmp_685;
  assign _mul_19_sink_stop = _tmp_685;
  reg _tmp_686;
  reg _tmp_687;
  reg _tmp_688;
  reg _tmp_689;
  reg _tmp_690;
  reg _tmp_691;
  reg _tmp_692;
  reg _tmp_693;
  reg _tmp_694;
  reg _tmp_695;
  assign _mul_19_sink_busy = _tmp_695;
  reg _tmp_696;
  assign _mul_19_busy = _mul_19_source_busy || _mul_19_sink_busy || _mul_19_busy_reg;
  reg _tmp_697;
  reg _tmp_698;
  reg _tmp_699;
  assign _mul_20_source_stop = _mul_20_stream_oready && 1'd0;
  reg _tmp_700;
  reg _tmp_701;
  reg _tmp_702;
  reg _tmp_703;
  reg _tmp_704;
  reg _tmp_705;
  reg _tmp_706;
  reg _tmp_707;
  reg _tmp_708;
  reg _tmp_709;
  assign _mul_20_sink_start = _tmp_709;
  reg _tmp_710;
  reg _tmp_711;
  reg _tmp_712;
  reg _tmp_713;
  reg _tmp_714;
  reg _tmp_715;
  reg _tmp_716;
  reg _tmp_717;
  reg _tmp_718;
  reg _tmp_719;
  assign _mul_20_sink_stop = _tmp_719;
  reg _tmp_720;
  reg _tmp_721;
  reg _tmp_722;
  reg _tmp_723;
  reg _tmp_724;
  reg _tmp_725;
  reg _tmp_726;
  reg _tmp_727;
  reg _tmp_728;
  reg _tmp_729;
  assign _mul_20_sink_busy = _tmp_729;
  reg _tmp_730;
  assign _mul_20_busy = _mul_20_source_busy || _mul_20_sink_busy || _mul_20_busy_reg;
  reg _tmp_731;
  reg _tmp_732;
  reg _tmp_733;
  assign _mul_21_source_stop = _mul_21_stream_oready && 1'd0;
  reg _tmp_734;
  reg _tmp_735;
  reg _tmp_736;
  reg _tmp_737;
  reg _tmp_738;
  reg _tmp_739;
  reg _tmp_740;
  reg _tmp_741;
  reg _tmp_742;
  reg _tmp_743;
  assign _mul_21_sink_start = _tmp_743;
  reg _tmp_744;
  reg _tmp_745;
  reg _tmp_746;
  reg _tmp_747;
  reg _tmp_748;
  reg _tmp_749;
  reg _tmp_750;
  reg _tmp_751;
  reg _tmp_752;
  reg _tmp_753;
  assign _mul_21_sink_stop = _tmp_753;
  reg _tmp_754;
  reg _tmp_755;
  reg _tmp_756;
  reg _tmp_757;
  reg _tmp_758;
  reg _tmp_759;
  reg _tmp_760;
  reg _tmp_761;
  reg _tmp_762;
  reg _tmp_763;
  assign _mul_21_sink_busy = _tmp_763;
  reg _tmp_764;
  assign _mul_21_busy = _mul_21_source_busy || _mul_21_sink_busy || _mul_21_busy_reg;
  reg _tmp_765;
  reg _tmp_766;
  reg _tmp_767;
  assign _mul_22_source_stop = _mul_22_stream_oready && 1'd0;
  reg _tmp_768;
  reg _tmp_769;
  reg _tmp_770;
  reg _tmp_771;
  reg _tmp_772;
  reg _tmp_773;
  reg _tmp_774;
  reg _tmp_775;
  reg _tmp_776;
  reg _tmp_777;
  assign _mul_22_sink_start = _tmp_777;
  reg _tmp_778;
  reg _tmp_779;
  reg _tmp_780;
  reg _tmp_781;
  reg _tmp_782;
  reg _tmp_783;
  reg _tmp_784;
  reg _tmp_785;
  reg _tmp_786;
  reg _tmp_787;
  assign _mul_22_sink_stop = _tmp_787;
  reg _tmp_788;
  reg _tmp_789;
  reg _tmp_790;
  reg _tmp_791;
  reg _tmp_792;
  reg _tmp_793;
  reg _tmp_794;
  reg _tmp_795;
  reg _tmp_796;
  reg _tmp_797;
  assign _mul_22_sink_busy = _tmp_797;
  reg _tmp_798;
  assign _mul_22_busy = _mul_22_source_busy || _mul_22_sink_busy || _mul_22_busy_reg;
  reg _tmp_799;
  reg _tmp_800;
  reg _tmp_801;
  assign _mul_23_source_stop = _mul_23_stream_oready && 1'd0;
  reg _tmp_802;
  reg _tmp_803;
  reg _tmp_804;
  reg _tmp_805;
  reg _tmp_806;
  reg _tmp_807;
  reg _tmp_808;
  reg _tmp_809;
  reg _tmp_810;
  reg _tmp_811;
  assign _mul_23_sink_start = _tmp_811;
  reg _tmp_812;
  reg _tmp_813;
  reg _tmp_814;
  reg _tmp_815;
  reg _tmp_816;
  reg _tmp_817;
  reg _tmp_818;
  reg _tmp_819;
  reg _tmp_820;
  reg _tmp_821;
  assign _mul_23_sink_stop = _tmp_821;
  reg _tmp_822;
  reg _tmp_823;
  reg _tmp_824;
  reg _tmp_825;
  reg _tmp_826;
  reg _tmp_827;
  reg _tmp_828;
  reg _tmp_829;
  reg _tmp_830;
  reg _tmp_831;
  assign _mul_23_sink_busy = _tmp_831;
  reg _tmp_832;
  assign _mul_23_busy = _mul_23_source_busy || _mul_23_sink_busy || _mul_23_busy_reg;
  reg _tmp_833;
  reg _tmp_834;
  reg _tmp_835;
  assign _mul_24_source_stop = _mul_24_stream_oready && 1'd0;
  reg _tmp_836;
  reg _tmp_837;
  reg _tmp_838;
  reg _tmp_839;
  reg _tmp_840;
  reg _tmp_841;
  reg _tmp_842;
  reg _tmp_843;
  reg _tmp_844;
  reg _tmp_845;
  assign _mul_24_sink_start = _tmp_845;
  reg _tmp_846;
  reg _tmp_847;
  reg _tmp_848;
  reg _tmp_849;
  reg _tmp_850;
  reg _tmp_851;
  reg _tmp_852;
  reg _tmp_853;
  reg _tmp_854;
  reg _tmp_855;
  assign _mul_24_sink_stop = _tmp_855;
  reg _tmp_856;
  reg _tmp_857;
  reg _tmp_858;
  reg _tmp_859;
  reg _tmp_860;
  reg _tmp_861;
  reg _tmp_862;
  reg _tmp_863;
  reg _tmp_864;
  reg _tmp_865;
  assign _mul_24_sink_busy = _tmp_865;
  reg _tmp_866;
  assign _mul_24_busy = _mul_24_source_busy || _mul_24_sink_busy || _mul_24_busy_reg;
  reg _tmp_867;
  reg _tmp_868;
  reg _tmp_869;
  assign _mul_25_source_stop = _mul_25_stream_oready && 1'd0;
  reg _tmp_870;
  reg _tmp_871;
  reg _tmp_872;
  reg _tmp_873;
  reg _tmp_874;
  reg _tmp_875;
  reg _tmp_876;
  reg _tmp_877;
  reg _tmp_878;
  reg _tmp_879;
  assign _mul_25_sink_start = _tmp_879;
  reg _tmp_880;
  reg _tmp_881;
  reg _tmp_882;
  reg _tmp_883;
  reg _tmp_884;
  reg _tmp_885;
  reg _tmp_886;
  reg _tmp_887;
  reg _tmp_888;
  reg _tmp_889;
  assign _mul_25_sink_stop = _tmp_889;
  reg _tmp_890;
  reg _tmp_891;
  reg _tmp_892;
  reg _tmp_893;
  reg _tmp_894;
  reg _tmp_895;
  reg _tmp_896;
  reg _tmp_897;
  reg _tmp_898;
  reg _tmp_899;
  assign _mul_25_sink_busy = _tmp_899;
  reg _tmp_900;
  assign _mul_25_busy = _mul_25_source_busy || _mul_25_sink_busy || _mul_25_busy_reg;
  reg _tmp_901;
  reg _tmp_902;
  reg _tmp_903;
  assign _mul_26_source_stop = _mul_26_stream_oready && 1'd0;
  reg _tmp_904;
  reg _tmp_905;
  reg _tmp_906;
  reg _tmp_907;
  reg _tmp_908;
  reg _tmp_909;
  reg _tmp_910;
  reg _tmp_911;
  reg _tmp_912;
  reg _tmp_913;
  assign _mul_26_sink_start = _tmp_913;
  reg _tmp_914;
  reg _tmp_915;
  reg _tmp_916;
  reg _tmp_917;
  reg _tmp_918;
  reg _tmp_919;
  reg _tmp_920;
  reg _tmp_921;
  reg _tmp_922;
  reg _tmp_923;
  assign _mul_26_sink_stop = _tmp_923;
  reg _tmp_924;
  reg _tmp_925;
  reg _tmp_926;
  reg _tmp_927;
  reg _tmp_928;
  reg _tmp_929;
  reg _tmp_930;
  reg _tmp_931;
  reg _tmp_932;
  reg _tmp_933;
  assign _mul_26_sink_busy = _tmp_933;
  reg _tmp_934;
  assign _mul_26_busy = _mul_26_source_busy || _mul_26_sink_busy || _mul_26_busy_reg;
  reg _tmp_935;
  reg _tmp_936;
  reg _tmp_937;
  assign _add_tree_16_source_stop = _add_tree_16_stream_oready && 1'd0;
  reg _tmp_938;
  reg _tmp_939;
  reg _tmp_940;
  reg _tmp_941;
  assign _add_tree_16_sink_start = _tmp_941;
  reg _tmp_942;
  reg _tmp_943;
  reg _tmp_944;
  reg _tmp_945;
  assign _add_tree_16_sink_stop = _tmp_945;
  reg _tmp_946;
  reg _tmp_947;
  reg _tmp_948;
  reg _tmp_949;
  assign _add_tree_16_sink_busy = _tmp_949;
  reg _tmp_950;
  assign _add_tree_16_busy = _add_tree_16_source_busy || _add_tree_16_sink_busy || _add_tree_16_busy_reg;
  reg _tmp_951;
  reg _tmp_952;
  reg _tmp_953;
  reg _tmp_954;
  reg _tmp_955;
  reg _tmp_956;
  reg _tmp_957;
  reg _tmp_958;
  reg _tmp_959;
  reg _tmp_960;
  assign _acc_14_source_stop = _acc_14_stream_oready && 1'd0;
  reg _tmp_961;
  reg _tmp_962;
  reg _tmp_963;
  reg _tmp_964;
  reg _tmp_965;
  reg _tmp_966;
  reg _tmp_967;
  assign _acc_14_sink_start = _tmp_967;
  reg _tmp_968;
  reg _tmp_969;
  reg _tmp_970;
  reg _tmp_971;
  reg _tmp_972;
  reg _tmp_973;
  reg _tmp_974;
  assign _acc_14_sink_stop = _tmp_974;
  reg _tmp_975;
  reg _tmp_976;
  reg _tmp_977;
  reg _tmp_978;
  reg _tmp_979;
  reg _tmp_980;
  reg _tmp_981;
  assign _acc_14_sink_busy = _tmp_981;
  reg _tmp_982;
  assign _acc_14_busy = _acc_14_source_busy || _acc_14_sink_busy || _acc_14_busy_reg;
  reg _tmp_983;
  reg _tmp_984;
  reg _tmp_985;
  assign _mul_rshift_round_clip_17_source_stop = _mul_rshift_round_clip_17_stream_oready && 1'd0;
  reg _tmp_986;
  reg _tmp_987;
  reg _tmp_988;
  reg _tmp_989;
  reg _tmp_990;
  reg _tmp_991;
  reg _tmp_992;
  reg _tmp_993;
  reg _tmp_994;
  reg _tmp_995;
  assign _mul_rshift_round_clip_17_sink_start = _tmp_995;
  reg _tmp_996;
  reg _tmp_997;
  reg _tmp_998;
  reg _tmp_999;
  reg _tmp_1000;
  reg _tmp_1001;
  reg _tmp_1002;
  reg _tmp_1003;
  reg _tmp_1004;
  reg _tmp_1005;
  assign _mul_rshift_round_clip_17_sink_stop = _tmp_1005;
  reg _tmp_1006;
  reg _tmp_1007;
  reg _tmp_1008;
  reg _tmp_1009;
  reg _tmp_1010;
  reg _tmp_1011;
  reg _tmp_1012;
  reg _tmp_1013;
  reg _tmp_1014;
  reg _tmp_1015;
  assign _mul_rshift_round_clip_17_sink_busy = _tmp_1015;
  reg _tmp_1016;
  assign _mul_rshift_round_clip_17_busy = _mul_rshift_round_clip_17_source_busy || _mul_rshift_round_clip_17_sink_busy || _mul_rshift_round_clip_17_busy_reg;
  reg _tmp_1017;
  reg _tmp_1018;
  reg _tmp_1019;
  reg _tmp_1020;
  reg _tmp_1021;
  reg _tmp_1022;
  reg [1-1:0] __variable_wdata_1553;
  assign stream_conv2d_4__reduce_reset_data = __variable_wdata_1553;
  reg _tmp_1023;
  reg _tmp_1024;
  reg _tmp_1025;
  reg _tmp_1026;
  assign _stream_conv2d_4_source_stop = _stream_conv2d_4_stream_oready && (_stream_conv2d_4_source_11_idle && _stream_conv2d_4_source_13_idle && _stream_conv2d_4_source_15_idle && _stream_conv2d_4_source_20_idle && _stream_conv2d_4_source_21_idle && _stream_conv2d_4_source_22_idle && _stream_conv2d_4_source_23_idle && _stream_conv2d_4_source_24_idle && _stream_conv2d_4_source_25_idle && _stream_conv2d_4_source_26_idle && _stream_conv2d_4_source_27_idle && _stream_conv2d_4_source_28_idle && _stream_conv2d_4_source_29_idle && _stream_conv2d_4_source_30_idle && _stream_conv2d_4_source_31_idle && _stream_conv2d_4_source_32_idle && _stream_conv2d_4_source_33_idle && _stream_conv2d_4_source_34_idle && _stream_conv2d_4_source_35_idle && _stream_conv2d_4_source_36_idle && _stream_conv2d_4_source_37_idle && _stream_conv2d_4_source_7_idle && _stream_conv2d_4_source_9_idle && (_stream_conv2d_4_fsm == 3));
  localparam _tmp_1027 = 1;
  wire [_tmp_1027-1:0] _tmp_1028;
  assign _tmp_1028 = _stream_conv2d_4_source_11_idle && _stream_conv2d_4_source_13_idle && _stream_conv2d_4_source_15_idle && _stream_conv2d_4_source_20_idle && _stream_conv2d_4_source_21_idle && _stream_conv2d_4_source_22_idle && _stream_conv2d_4_source_23_idle && _stream_conv2d_4_source_24_idle && _stream_conv2d_4_source_25_idle && _stream_conv2d_4_source_26_idle && _stream_conv2d_4_source_27_idle && _stream_conv2d_4_source_28_idle && _stream_conv2d_4_source_29_idle && _stream_conv2d_4_source_30_idle && _stream_conv2d_4_source_31_idle && _stream_conv2d_4_source_32_idle && _stream_conv2d_4_source_33_idle && _stream_conv2d_4_source_34_idle && _stream_conv2d_4_source_35_idle && _stream_conv2d_4_source_36_idle && _stream_conv2d_4_source_37_idle && _stream_conv2d_4_source_7_idle && _stream_conv2d_4_source_9_idle && (_stream_conv2d_4_fsm == 3);
  reg [_tmp_1027-1:0] _tmp_1029;
  localparam _tmp_1030 = 1;
  wire [_tmp_1030-1:0] _tmp_1031;
  assign _tmp_1031 = _stream_conv2d_4_source_11_idle && _stream_conv2d_4_source_13_idle && _stream_conv2d_4_source_15_idle && _stream_conv2d_4_source_20_idle && _stream_conv2d_4_source_21_idle && _stream_conv2d_4_source_22_idle && _stream_conv2d_4_source_23_idle && _stream_conv2d_4_source_24_idle && _stream_conv2d_4_source_25_idle && _stream_conv2d_4_source_26_idle && _stream_conv2d_4_source_27_idle && _stream_conv2d_4_source_28_idle && _stream_conv2d_4_source_29_idle && _stream_conv2d_4_source_30_idle && _stream_conv2d_4_source_31_idle && _stream_conv2d_4_source_32_idle && _stream_conv2d_4_source_33_idle && _stream_conv2d_4_source_34_idle && _stream_conv2d_4_source_35_idle && _stream_conv2d_4_source_36_idle && _stream_conv2d_4_source_37_idle && _stream_conv2d_4_source_7_idle && _stream_conv2d_4_source_9_idle && (_stream_conv2d_4_fsm == 3);
  reg [_tmp_1030-1:0] _tmp_1032;
  reg _tmp_1033;
  reg _tmp_1034;
  reg _tmp_1035;
  reg _tmp_1036;
  reg _tmp_1037;
  reg _tmp_1038;
  reg _tmp_1039;
  reg _tmp_1040;
  reg _tmp_1041;
  reg _tmp_1042;
  reg _tmp_1043;
  reg _tmp_1044;
  reg _tmp_1045;
  reg _tmp_1046;
  reg _tmp_1047;
  reg _tmp_1048;
  reg _tmp_1049;
  reg _tmp_1050;
  reg _tmp_1051;
  reg _tmp_1052;
  reg _tmp_1053;
  reg _tmp_1054;
  reg _tmp_1055;
  reg _tmp_1056;
  reg _tmp_1057;
  reg _tmp_1058;
  reg _tmp_1059;
  reg _tmp_1060;
  reg _tmp_1061;
  reg _tmp_1062;
  reg _tmp_1063;
  reg _tmp_1064;
  reg _tmp_1065;
  assign _stream_conv2d_4_sink_start = _tmp_1065;
  reg _tmp_1066;
  reg _tmp_1067;
  reg _tmp_1068;
  reg _tmp_1069;
  reg _tmp_1070;
  reg _tmp_1071;
  reg _tmp_1072;
  reg _tmp_1073;
  reg _tmp_1074;
  reg _tmp_1075;
  reg _tmp_1076;
  reg _tmp_1077;
  reg _tmp_1078;
  reg _tmp_1079;
  reg _tmp_1080;
  reg _tmp_1081;
  reg _tmp_1082;
  reg _tmp_1083;
  reg _tmp_1084;
  reg _tmp_1085;
  reg _tmp_1086;
  reg _tmp_1087;
  reg _tmp_1088;
  reg _tmp_1089;
  reg _tmp_1090;
  reg _tmp_1091;
  reg _tmp_1092;
  reg _tmp_1093;
  reg _tmp_1094;
  reg _tmp_1095;
  reg _tmp_1096;
  reg _tmp_1097;
  reg _tmp_1098;
  assign _stream_conv2d_4_sink_stop = _tmp_1098;
  reg _tmp_1099;
  reg _tmp_1100;
  reg _tmp_1101;
  reg _tmp_1102;
  reg _tmp_1103;
  reg _tmp_1104;
  reg _tmp_1105;
  reg _tmp_1106;
  reg _tmp_1107;
  reg _tmp_1108;
  reg _tmp_1109;
  reg _tmp_1110;
  reg _tmp_1111;
  reg _tmp_1112;
  reg _tmp_1113;
  reg _tmp_1114;
  reg _tmp_1115;
  reg _tmp_1116;
  reg _tmp_1117;
  reg _tmp_1118;
  reg _tmp_1119;
  reg _tmp_1120;
  reg _tmp_1121;
  reg _tmp_1122;
  reg _tmp_1123;
  reg _tmp_1124;
  reg _tmp_1125;
  reg _tmp_1126;
  reg _tmp_1127;
  reg _tmp_1128;
  reg _tmp_1129;
  reg _tmp_1130;
  reg _tmp_1131;
  assign _stream_conv2d_4_sink_busy = _tmp_1131;
  reg _tmp_1132;
  assign _stream_conv2d_4_busy = _stream_conv2d_4_source_busy || _stream_conv2d_4_sink_busy || _stream_conv2d_4_busy_reg;
  wire conv2d_4_dma_out_mask_0;
  assign conv2d_4_dma_out_mask_0 = conv2d_4_out_row_count + 0 >= cparam_conv2d_4_out_num_row;
  wire [32-1:0] _dma_write_packed_high_local_size_1133;
  assign _dma_write_packed_high_local_size_1133 = conv2d_4_next_out_write_size >> 1;
  wire [1-1:0] _dma_write_packed_low_local_size_1134;
  assign _dma_write_packed_low_local_size_1134 = conv2d_4_next_out_write_size & { 1{ 1'd1 } };
  wire [32-1:0] _dma_write_packed_local_packed_size_1135;
  assign _dma_write_packed_local_packed_size_1135 = (_dma_write_packed_low_local_size_1134 > 0)? _dma_write_packed_high_local_size_1133 + 1 : _dma_write_packed_high_local_size_1133;
  wire [32-1:0] mask_addr_shifted_1136;
  assign mask_addr_shifted_1136 = conv2d_4_objaddr + (conv2d_4_out_base_offset + cparam_conv2d_4_out_offset_values_0) + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_1137;
  assign mask_addr_masked_1137 = mask_addr_shifted_1136 << 2;
  reg [32-1:0] _maxi_write_req_fsm;
  localparam _maxi_write_req_fsm_init = 0;
  reg [33-1:0] _maxi_write_cur_global_size;
  reg _maxi_write_cont;
  wire [8-1:0] pack_write_req_op_sel_1138;
  wire [32-1:0] pack_write_req_local_addr_1139;
  wire [32-1:0] pack_write_req_local_stride_1140;
  wire [33-1:0] pack_write_req_size_1141;
  wire [32-1:0] pack_write_req_local_blocksize_1142;
  assign pack_write_req_op_sel_1138 = _maxi_write_op_sel;
  assign pack_write_req_local_addr_1139 = _maxi_write_local_addr;
  assign pack_write_req_local_stride_1140 = _maxi_write_local_stride;
  assign pack_write_req_size_1141 = _maxi_write_local_size;
  assign pack_write_req_local_blocksize_1142 = _maxi_write_local_blocksize;
  wire [137-1:0] pack_write_req_packed_1143;
  assign pack_write_req_packed_1143 = { pack_write_req_op_sel_1138, pack_write_req_local_addr_1139, pack_write_req_local_stride_1140, pack_write_req_size_1141, pack_write_req_local_blocksize_1142 };
  localparam _tmp_1144 = 1;
  wire [_tmp_1144-1:0] _tmp_1145;
  assign _tmp_1145 = !_maxi_write_req_fifo_almost_full;
  reg [_tmp_1144-1:0] __tmp_1145_1;
  wire [32-1:0] mask_addr_shifted_1146;
  assign mask_addr_shifted_1146 = _maxi_write_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_1147;
  assign mask_addr_masked_1147 = mask_addr_shifted_1146 << 2;
  wire [32-1:0] mask_addr_shifted_1148;
  assign mask_addr_shifted_1148 = _maxi_write_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_1149;
  assign mask_addr_masked_1149 = mask_addr_shifted_1148 << 2;
  wire [32-1:0] mask_addr_shifted_1150;
  assign mask_addr_shifted_1150 = _maxi_write_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_1151;
  assign mask_addr_masked_1151 = mask_addr_shifted_1150 << 2;
  wire [32-1:0] mask_addr_shifted_1152;
  assign mask_addr_shifted_1152 = _maxi_write_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_1153;
  assign mask_addr_masked_1153 = mask_addr_shifted_1152 << 2;
  wire [32-1:0] mask_addr_shifted_1154;
  assign mask_addr_shifted_1154 = _maxi_write_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_1155;
  assign mask_addr_masked_1155 = mask_addr_shifted_1154 << 2;
  wire [32-1:0] mask_addr_shifted_1156;
  assign mask_addr_shifted_1156 = _maxi_write_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_1157;
  assign mask_addr_masked_1157 = mask_addr_shifted_1156 << 2;
  wire [8-1:0] pack_write_req_op_sel_1158;
  wire [32-1:0] pack_write_req_local_addr_1159;
  wire [32-1:0] pack_write_req_local_stride_1160;
  wire [33-1:0] pack_write_req_size_1161;
  wire [32-1:0] pack_write_req_local_blocksize_1162;
  assign pack_write_req_op_sel_1158 = _maxi_write_op_sel;
  assign pack_write_req_local_addr_1159 = _maxi_write_local_addr;
  assign pack_write_req_local_stride_1160 = _maxi_write_local_stride;
  assign pack_write_req_size_1161 = _maxi_write_cur_global_size;
  assign pack_write_req_local_blocksize_1162 = _maxi_write_local_blocksize;
  wire [137-1:0] pack_write_req_packed_1163;
  assign pack_write_req_packed_1163 = { pack_write_req_op_sel_1158, pack_write_req_local_addr_1159, pack_write_req_local_stride_1160, pack_write_req_size_1161, pack_write_req_local_blocksize_1162 };
  assign _maxi_write_req_fifo_wdata = ((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (maxi_awready || !maxi_awvalid) && (_maxi_outstanding_wcount < 6))? pack_write_req_packed_1163 : 
                                      ((_maxi_write_req_fsm == 0) && _maxi_write_start && !_maxi_write_req_fifo_almost_full)? pack_write_req_packed_1143 : 'hx;
  assign _maxi_write_req_fifo_enq = ((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (maxi_awready || !maxi_awvalid) && (_maxi_outstanding_wcount < 6))? (_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (maxi_awready || !maxi_awvalid) && (_maxi_outstanding_wcount < 6) && !_maxi_write_req_fifo_almost_full : 
                                    ((_maxi_write_req_fsm == 0) && _maxi_write_start && !_maxi_write_req_fifo_almost_full)? (_maxi_write_req_fsm == 0) && _maxi_write_start && !_maxi_write_req_fifo_almost_full && !_maxi_write_req_fifo_almost_full : 0;
  localparam _tmp_1164 = 1;
  wire [_tmp_1164-1:0] _tmp_1165;
  assign _tmp_1165 = !_maxi_write_req_fifo_almost_full;
  reg [_tmp_1164-1:0] __tmp_1165_1;
  reg _maxi_waddr_cond_0_1;
  reg [32-1:0] _maxi_write_data_fsm;
  localparam _maxi_write_data_fsm_init = 0;
  reg [32-1:0] read_burst_packed_fsm_55;
  localparam read_burst_packed_fsm_55_init = 0;
  reg [9-1:0] read_burst_packed_addr_1166;
  reg [9-1:0] read_burst_packed_stride_1167;
  reg [33-1:0] read_burst_packed_length_1168;
  reg read_burst_packed_rvalid_1169;
  reg read_burst_packed_rlast_1170;
  wire [8-1:0] read_burst_packed_ram_addr_1171;
  assign read_burst_packed_ram_addr_1171 = read_burst_packed_addr_1166 >> 1;
  assign ram_w16_l512_id20_0_1_addr = ((read_burst_packed_fsm_55 == 1) && (!read_burst_packed_rvalid_1169 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? read_burst_packed_ram_addr_1171 : 'hx;
  assign ram_w16_l512_id20_0_1_enable = ((read_burst_packed_fsm_55 == 1) && (!read_burst_packed_rvalid_1169 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? 1'd1 : 0;
  localparam _tmp_1172 = 1;
  wire [_tmp_1172-1:0] _tmp_1173;
  assign _tmp_1173 = (read_burst_packed_fsm_55 == 1) && (!read_burst_packed_rvalid_1169 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0));
  reg [_tmp_1172-1:0] __tmp_1173_1;
  wire [16-1:0] read_burst_packed_ram_rdata_1174;
  assign read_burst_packed_ram_rdata_1174 = ram_w16_l512_id20_0_1_rdata;
  wire [8-1:0] read_burst_packed_ram_addr_1175;
  assign read_burst_packed_ram_addr_1175 = read_burst_packed_addr_1166 >> 1;
  assign ram_w16_l512_id20_1_1_addr = ((read_burst_packed_fsm_55 == 1) && (!read_burst_packed_rvalid_1169 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? read_burst_packed_ram_addr_1175 : 'hx;
  assign ram_w16_l512_id20_1_1_enable = ((read_burst_packed_fsm_55 == 1) && (!read_burst_packed_rvalid_1169 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? 1'd1 : 0;
  localparam _tmp_1176 = 1;
  wire [_tmp_1176-1:0] _tmp_1177;
  assign _tmp_1177 = (read_burst_packed_fsm_55 == 1) && (!read_burst_packed_rvalid_1169 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0));
  reg [_tmp_1176-1:0] __tmp_1177_1;
  wire [16-1:0] read_burst_packed_ram_rdata_1178;
  assign read_burst_packed_ram_rdata_1178 = ram_w16_l512_id20_1_1_rdata;
  wire [32-1:0] read_burst_packed_rdata_1179;
  assign read_burst_packed_rdata_1179 = { read_burst_packed_ram_rdata_1178, read_burst_packed_ram_rdata_1174 };
  reg _maxi_wdata_cond_0_1;
  wire conv2d_4_update_filter;
  assign conv2d_4_update_filter = (cparam_conv2d_4_data_stationary == 0) && (conv2d_4_row_count >= cparam_conv2d_4_max_row_count) && (conv2d_4_bat_count >= cparam_conv2d_4_max_bat_count) || (cparam_conv2d_4_data_stationary == 1) && !cparam_conv2d_4_keep_filter;
  wire conv2d_4_update_act;
  assign conv2d_4_update_act = (cparam_conv2d_4_data_stationary == 1) && (conv2d_4_och_count >= cparam_conv2d_4_max_och_count) || (cparam_conv2d_4_data_stationary == 0);
  wire conv2d_4_mux_next_dma_flag_0;
  assign conv2d_4_mux_next_dma_flag_0 = (conv2d_4_row_select == 0)? (conv2d_4_row_count >= cparam_conv2d_4_max_row_count)? 1 : cparam_conv2d_4_dma_flag_conds_0 : 
                                        (conv2d_4_row_select == 1)? (conv2d_4_row_count >= cparam_conv2d_4_max_row_count)? 1 : cparam_conv2d_4_dma_flag_conds_2 : 
                                        (conv2d_4_row_select == 2)? (conv2d_4_row_count >= cparam_conv2d_4_max_row_count)? 1 : cparam_conv2d_4_dma_flag_conds_1 : 1'd0;
  wire conv2d_4_mux_next_dma_flag_1;
  assign conv2d_4_mux_next_dma_flag_1 = (conv2d_4_row_select == 0)? (conv2d_4_row_count >= cparam_conv2d_4_max_row_count)? 1 : cparam_conv2d_4_dma_flag_conds_1 : 
                                        (conv2d_4_row_select == 1)? (conv2d_4_row_count >= cparam_conv2d_4_max_row_count)? 1 : cparam_conv2d_4_dma_flag_conds_0 : 
                                        (conv2d_4_row_select == 2)? (conv2d_4_row_count >= cparam_conv2d_4_max_row_count)? 1 : cparam_conv2d_4_dma_flag_conds_2 : 1'd0;
  wire conv2d_4_mux_next_dma_flag_2;
  assign conv2d_4_mux_next_dma_flag_2 = (conv2d_4_row_select == 0)? (conv2d_4_row_count >= cparam_conv2d_4_max_row_count)? 1 : cparam_conv2d_4_dma_flag_conds_2 : 
                                        (conv2d_4_row_select == 1)? (conv2d_4_row_count >= cparam_conv2d_4_max_row_count)? 1 : cparam_conv2d_4_dma_flag_conds_1 : 
                                        (conv2d_4_row_select == 2)? (conv2d_4_row_count >= cparam_conv2d_4_max_row_count)? 1 : cparam_conv2d_4_dma_flag_conds_0 : 1'd0;
  reg [32-1:0] max_pool_serial_6_objaddr;
  reg [32-1:0] max_pool_serial_6_arg_objaddr_0;
  reg [32-1:0] control_max_pool_serial_6;
  localparam control_max_pool_serial_6_init = 0;
  reg _control_max_pool_serial_6_called;
  wire signed [32-1:0] max_pool_serial_6_act_base_offset;
  reg signed [32-1:0] max_pool_serial_6_act_base_offset_row;
  reg signed [32-1:0] max_pool_serial_6_act_base_offset_bat;
  assign max_pool_serial_6_act_base_offset = max_pool_serial_6_act_base_offset_row + max_pool_serial_6_act_base_offset_bat;
  wire signed [32-1:0] max_pool_serial_6_out_base_offset;
  reg signed [32-1:0] max_pool_serial_6_out_base_offset_row;
  reg signed [32-1:0] max_pool_serial_6_out_base_offset_bat;
  assign max_pool_serial_6_out_base_offset = max_pool_serial_6_out_base_offset_row + max_pool_serial_6_out_base_offset_bat;
  reg [32-1:0] max_pool_serial_6_col_count;
  reg [32-1:0] max_pool_serial_6_row_count;
  reg [32-1:0] max_pool_serial_6_bat_count;
  reg [32-1:0] max_pool_serial_6_prev_row_count;
  reg [32-1:0] max_pool_serial_6_prev_bat_count;
  reg [32-1:0] max_pool_serial_6_stream_act_local;
  reg [32-1:0] max_pool_serial_6_stream_out_local;
  reg max_pool_serial_6_act_page;
  reg [32-1:0] max_pool_serial_6_act_page_comp_offset;
  reg [32-1:0] max_pool_serial_6_act_page_dma_offset;
  reg max_pool_serial_6_out_page;
  reg [32-1:0] max_pool_serial_6_out_page_comp_offset;
  reg [32-1:0] max_pool_serial_6_out_page_dma_offset;
  reg max_pool_serial_6_skip_read_act;
  reg max_pool_serial_6_skip_comp;
  reg max_pool_serial_6_skip_write_out;
  reg [32-1:0] max_pool_serial_6_comp_count;
  reg [32-1:0] max_pool_serial_6_out_count;
  wire max_pool_serial_6_dma_pad_mask_0;
  assign max_pool_serial_6_dma_pad_mask_0 = (max_pool_serial_6_row_count + 0 < cparam_max_pool_serial_6_pad_row_top) || (max_pool_serial_6_row_count + 0 >= cparam_max_pool_serial_6_act_num_row + cparam_max_pool_serial_6_pad_row_top);
  wire max_pool_serial_6_dma_pad_mask_1;
  assign max_pool_serial_6_dma_pad_mask_1 = (max_pool_serial_6_row_count + 1 < cparam_max_pool_serial_6_pad_row_top) || (max_pool_serial_6_row_count + 1 >= cparam_max_pool_serial_6_act_num_row + cparam_max_pool_serial_6_pad_row_top);
  wire [10-1:0] _dma_read_packed_high_local_size_1180;
  assign _dma_read_packed_high_local_size_1180 = cparam_max_pool_serial_6_act_read_size >> 1;
  wire [1-1:0] _dma_read_packed_low_local_size_1181;
  assign _dma_read_packed_low_local_size_1181 = cparam_max_pool_serial_6_act_read_size & { 1{ 1'd1 } };
  wire [10-1:0] _dma_read_packed_local_packed_size_1182;
  assign _dma_read_packed_local_packed_size_1182 = (_dma_read_packed_low_local_size_1181 > 0)? _dma_read_packed_high_local_size_1180 + 1 : _dma_read_packed_high_local_size_1180;
  wire [32-1:0] mask_addr_shifted_1183;
  assign mask_addr_shifted_1183 = max_pool_serial_6_arg_objaddr_0 + (max_pool_serial_6_act_base_offset + cparam_max_pool_serial_6_act_offset_values_0) + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_1184;
  assign mask_addr_masked_1184 = mask_addr_shifted_1183 << 2;
  reg [32-1:0] write_burst_packed_fsm_56;
  localparam write_burst_packed_fsm_56_init = 0;
  reg [15-1:0] write_burst_packed_addr_1185;
  reg [15-1:0] write_burst_packed_stride_1186;
  reg [33-1:0] write_burst_packed_length_1187;
  reg write_burst_packed_done_1188;
  wire [14-1:0] write_burst_packed_ram_addr_1189;
  assign write_burst_packed_ram_addr_1189 = write_burst_packed_addr_1185 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_1190;
  assign write_burst_packed_ram_wdata_1190 = _maxi_rdata_sb_0 >> 0;
  assign ram_w16_l32768_id0_0_1_addr = ((write_burst_packed_fsm_56 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_addr_1189 : 'hx;
  assign ram_w16_l32768_id0_0_1_wdata = ((write_burst_packed_fsm_56 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_wdata_1190 : 'hx;
  assign ram_w16_l32768_id0_0_1_wenable = ((write_burst_packed_fsm_56 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  assign ram_w16_l32768_id0_0_1_enable = ((write_burst_packed_fsm_56 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  wire [14-1:0] write_burst_packed_ram_addr_1191;
  assign write_burst_packed_ram_addr_1191 = write_burst_packed_addr_1185 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_1192;
  assign write_burst_packed_ram_wdata_1192 = _maxi_rdata_sb_0 >> 16;
  assign ram_w16_l32768_id0_1_1_addr = ((write_burst_packed_fsm_56 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_addr_1191 : 'hx;
  assign ram_w16_l32768_id0_1_1_wdata = ((write_burst_packed_fsm_56 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_wdata_1192 : 'hx;
  assign ram_w16_l32768_id0_1_1_wenable = ((write_burst_packed_fsm_56 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  assign ram_w16_l32768_id0_1_1_enable = ((write_burst_packed_fsm_56 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  wire [10-1:0] _dma_read_packed_high_local_size_1193;
  assign _dma_read_packed_high_local_size_1193 = cparam_max_pool_serial_6_act_read_size >> 1;
  wire [1-1:0] _dma_read_packed_low_local_size_1194;
  assign _dma_read_packed_low_local_size_1194 = cparam_max_pool_serial_6_act_read_size & { 1{ 1'd1 } };
  wire [10-1:0] _dma_read_packed_local_packed_size_1195;
  assign _dma_read_packed_local_packed_size_1195 = (_dma_read_packed_low_local_size_1194 > 0)? _dma_read_packed_high_local_size_1193 + 1 : _dma_read_packed_high_local_size_1193;
  wire [32-1:0] mask_addr_shifted_1196;
  assign mask_addr_shifted_1196 = max_pool_serial_6_arg_objaddr_0 + (max_pool_serial_6_act_base_offset + cparam_max_pool_serial_6_act_offset_values_1) + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_1197;
  assign mask_addr_masked_1197 = mask_addr_shifted_1196 << 2;
  reg [32-1:0] max_pool_serial_6_comp_fsm;
  localparam max_pool_serial_6_comp_fsm_init = 0;
  reg [32-1:0] max_pool_serial_6_act_page_comp_offset_buf;
  reg [32-1:0] max_pool_serial_6_out_page_comp_offset_buf;
  reg [32-1:0] max_pool_serial_6_row_count_buf;
  wire max_pool_serial_6_stream_pad_mask_0_0;
  assign max_pool_serial_6_stream_pad_mask_0_0 = (max_pool_serial_6_col_count + 0 < cparam_max_pool_serial_6_pad_col_left) || (max_pool_serial_6_col_count + 0 >= cparam_max_pool_serial_6_act_num_col + cparam_max_pool_serial_6_pad_col_left) || (max_pool_serial_6_row_count_buf + 0 < cparam_max_pool_serial_6_pad_row_top) || (max_pool_serial_6_row_count_buf + 0 >= cparam_max_pool_serial_6_act_num_row + cparam_max_pool_serial_6_pad_row_top);
  wire max_pool_serial_6_stream_pad_mask_0_1;
  assign max_pool_serial_6_stream_pad_mask_0_1 = (max_pool_serial_6_col_count + 1 < cparam_max_pool_serial_6_pad_col_left) || (max_pool_serial_6_col_count + 1 >= cparam_max_pool_serial_6_act_num_col + cparam_max_pool_serial_6_pad_col_left) || (max_pool_serial_6_row_count_buf + 0 < cparam_max_pool_serial_6_pad_row_top) || (max_pool_serial_6_row_count_buf + 0 >= cparam_max_pool_serial_6_act_num_row + cparam_max_pool_serial_6_pad_row_top);
  wire max_pool_serial_6_stream_pad_mask_1_0;
  assign max_pool_serial_6_stream_pad_mask_1_0 = (max_pool_serial_6_col_count + 0 < cparam_max_pool_serial_6_pad_col_left) || (max_pool_serial_6_col_count + 0 >= cparam_max_pool_serial_6_act_num_col + cparam_max_pool_serial_6_pad_col_left) || (max_pool_serial_6_row_count_buf + 1 < cparam_max_pool_serial_6_pad_row_top) || (max_pool_serial_6_row_count_buf + 1 >= cparam_max_pool_serial_6_act_num_row + cparam_max_pool_serial_6_pad_row_top);
  wire max_pool_serial_6_stream_pad_mask_1_1;
  assign max_pool_serial_6_stream_pad_mask_1_1 = (max_pool_serial_6_col_count + 1 < cparam_max_pool_serial_6_pad_col_left) || (max_pool_serial_6_col_count + 1 >= cparam_max_pool_serial_6_act_num_col + cparam_max_pool_serial_6_pad_col_left) || (max_pool_serial_6_row_count_buf + 1 < cparam_max_pool_serial_6_pad_row_top) || (max_pool_serial_6_row_count_buf + 1 >= cparam_max_pool_serial_6_act_num_row + cparam_max_pool_serial_6_pad_row_top);
  reg [4-1:0] max_pool_serial_6_stream_pad_masks;
  wire [3-1:0] stream_max_pool_serial_6_parameter_0_data;
  wire [16-1:0] stream_max_pool_serial_6_source_1_data;
  wire [4-1:0] stream_max_pool_serial_6_parameter_2_data;
  wire [1-1:0] stream_max_pool_serial_6__reduce_reset_data;
  reg __stream_max_pool_serial_6_stream_ivalid_1;
  reg __stream_max_pool_serial_6_stream_ivalid_2;
  reg __stream_max_pool_serial_6_stream_ivalid_3;
  reg __stream_max_pool_serial_6_stream_ivalid_4;
  reg __stream_max_pool_serial_6_stream_ivalid_5;
  reg [32-1:0] _counter_data_2141;
  reg [32-1:0] _counter_count_2141;
  wire _counter_reset_cond_2141;
  assign _counter_reset_cond_2141 = stream_max_pool_serial_6__reduce_reset_data;
  wire [32-1:0] _counter_current_count_2141;
  assign _counter_current_count_2141 = (_counter_reset_cond_2141)? 1'sd0 : _counter_count_2141;
  wire [16-1:0] _reinterpretcast_src_2149;
  assign _reinterpretcast_src_2149 = stream_max_pool_serial_6_source_1_data;
  wire signed [16-1:0] _reinterpretcast_data_2149;
  assign _reinterpretcast_data_2149 = _reinterpretcast_src_2149;
  reg [4-1:0] __delay_data_2394__variable_2139;
  reg signed [16-1:0] __delay_data_2395_reinterpretcast_2149;
  reg [1-1:0] __delay_data_2397__variable_2140;
  reg [3-1:0] __delay_data_2400__variable_2137;
  reg [1-1:0] _pointer_data_2144;
  reg signed [16-1:0] __delay_data_2396__delay_2395_reinterpretcast_2149;
  reg [1-1:0] __delay_data_2398__delay_2397__variable_2140;
  reg [3-1:0] __delay_data_2401__delay_2400__variable_2137;
  reg signed [17-1:0] _cond_data_2151;
  reg [1-1:0] __delay_data_2399__delay_2398__delay_2397__variable_2140;
  reg [3-1:0] __delay_data_2402__delay_2401__delay_2400__variable_2137;
  reg [1-1:0] __variable_wdata_1543;
  assign _reduce_max_27__reduce_reset_data = __variable_wdata_1543;
  reg signed [16-1:0] __variable_wdata_1541;
  assign _reduce_max_27_x_data = __variable_wdata_1541;
  reg [32-1:0] __variable_wdata_1542;
  assign _reduce_max_27_size_data = __variable_wdata_1542;
  assign __reduce_max_27_is_root = ((_stream_max_pool_serial_6_busy)? 0 : 1) && 1;
  assign __reduce_max_27_stream_oready = ((_stream_max_pool_serial_6_busy)? _stream_max_pool_serial_6_stream_oready : 1) && __reduce_max_27_stream_internal_oready;
  assign _stream_max_pool_serial_6_stream_internal_oready = ((_stream_max_pool_serial_6_busy)? __reduce_max_27_stream_internal_oready : 1) && 1;
  wire signed [16-1:0] __substreamoutput_data_2153;
  assign __substreamoutput_data_2153 = _reduce_max_27_data_data;
  wire [1-1:0] __substreamoutput_data_2154;
  assign __substreamoutput_data_2154 = _reduce_max_27_valid_data;
  wire signed [16-1:0] _reinterpretcast_src_2155;
  assign _reinterpretcast_src_2155 = __substreamoutput_data_2153;
  wire signed [16-1:0] _reinterpretcast_data_2155;
  assign _reinterpretcast_data_2155 = _reinterpretcast_src_2155;
  wire [1-1:0] stream_max_pool_serial_6_sink_6_data;
  assign stream_max_pool_serial_6_sink_6_data = __substreamoutput_data_2154;
  wire signed [16-1:0] stream_max_pool_serial_6_sink_5_data;
  assign stream_max_pool_serial_6_sink_5_data = _reinterpretcast_data_2155;
  wire _set_flag_1198;
  assign _set_flag_1198 = max_pool_serial_6_comp_fsm == 4;
  reg [3-1:0] __variable_wdata_2137;
  assign stream_max_pool_serial_6_parameter_0_data = __variable_wdata_2137;
  wire _set_flag_1199;
  assign _set_flag_1199 = max_pool_serial_6_comp_fsm == 4;
  reg [4-1:0] __variable_wdata_2139;
  assign stream_max_pool_serial_6_parameter_2_data = __variable_wdata_2139;
  reg [32-1:0] _source_stream_max_pool_serial_6_source_1_pat_cur_offset_0;
  reg [32-1:0] _source_stream_max_pool_serial_6_source_1_pat_cur_offset_1;
  reg [32-1:0] _source_stream_max_pool_serial_6_source_1_pat_cur_offset_2;
  reg [32-1:0] _source_stream_max_pool_serial_6_source_1_pat_cur_offset_3;
  reg [33-1:0] _source_stream_max_pool_serial_6_source_1_pat_size_0;
  reg [33-1:0] _source_stream_max_pool_serial_6_source_1_pat_size_1;
  reg [33-1:0] _source_stream_max_pool_serial_6_source_1_pat_size_2;
  reg [33-1:0] _source_stream_max_pool_serial_6_source_1_pat_size_3;
  reg [32-1:0] _source_stream_max_pool_serial_6_source_1_pat_stride_0;
  reg [32-1:0] _source_stream_max_pool_serial_6_source_1_pat_stride_1;
  reg [32-1:0] _source_stream_max_pool_serial_6_source_1_pat_stride_2;
  reg [32-1:0] _source_stream_max_pool_serial_6_source_1_pat_stride_3;
  reg [33-1:0] _source_stream_max_pool_serial_6_source_1_pat_count_0;
  reg [33-1:0] _source_stream_max_pool_serial_6_source_1_pat_count_1;
  reg [33-1:0] _source_stream_max_pool_serial_6_source_1_pat_count_2;
  reg [33-1:0] _source_stream_max_pool_serial_6_source_1_pat_count_3;
  reg [33-1:0] _source_stream_max_pool_serial_6_source_1_pat_size_buf_0;
  reg [33-1:0] _source_stream_max_pool_serial_6_source_1_pat_size_buf_1;
  reg [33-1:0] _source_stream_max_pool_serial_6_source_1_pat_size_buf_2;
  reg [33-1:0] _source_stream_max_pool_serial_6_source_1_pat_size_buf_3;
  reg [32-1:0] _source_stream_max_pool_serial_6_source_1_pat_stride_buf_0;
  reg [32-1:0] _source_stream_max_pool_serial_6_source_1_pat_stride_buf_1;
  reg [32-1:0] _source_stream_max_pool_serial_6_source_1_pat_stride_buf_2;
  reg [32-1:0] _source_stream_max_pool_serial_6_source_1_pat_stride_buf_3;
  wire _set_flag_1200;
  assign _set_flag_1200 = max_pool_serial_6_comp_fsm == 4;
  wire [1-1:0] read_rtl_bank_1201;
  assign read_rtl_bank_1201 = _stream_max_pool_serial_6_source_1_source_ram_raddr;
  reg [1-1:0] _tmp_1202;
  localparam _tmp_1203 = 1;
  wire [_tmp_1203-1:0] _tmp_1204;
  assign _tmp_1204 = _stream_max_pool_serial_6_stream_oready && _stream_max_pool_serial_6_source_1_source_ram_renable && (_stream_max_pool_serial_6_source_1_source_sel == 1);
  reg [_tmp_1203-1:0] __tmp_1204_1;
  localparam _tmp_1205 = 1;
  wire [_tmp_1205-1:0] _tmp_1206;
  assign _tmp_1206 = _stream_max_pool_serial_6_stream_oready && _stream_max_pool_serial_6_source_1_source_ram_renable && (_stream_max_pool_serial_6_source_1_source_sel == 1);
  reg [_tmp_1205-1:0] __tmp_1206_1;
  wire signed [16-1:0] read_rtl_rdata_1207;
  wire read_rtl_rvalid_1208;
  assign read_rtl_rdata_1207 = (_tmp_1202 == 0)? ram_w16_l32768_id0_0_0_rdata : 
                               (_tmp_1202 == 1)? ram_w16_l32768_id0_1_0_rdata : 0;
  assign read_rtl_rvalid_1208 = __tmp_1204_1;
  assign _stream_max_pool_serial_6_source_1_source_ram_rdata = (_stream_max_pool_serial_6_source_1_source_sel == 1)? read_rtl_rdata_1207 : 'hx;
  reg [16-1:0] __variable_wdata_2138;
  assign stream_max_pool_serial_6_source_1_data = __variable_wdata_2138;
  reg [32-1:0] _stream_max_pool_serial_6_source_1_source_pat_fsm_0;
  localparam _stream_max_pool_serial_6_source_1_source_pat_fsm_0_init = 0;
  wire [32-1:0] _stream_max_pool_serial_6_source_1_source_pat_all_offset;
  assign _stream_max_pool_serial_6_source_1_source_pat_all_offset = _stream_max_pool_serial_6_source_1_source_offset_buf + _source_stream_max_pool_serial_6_source_1_pat_cur_offset_0 + _source_stream_max_pool_serial_6_source_1_pat_cur_offset_1 + _source_stream_max_pool_serial_6_source_1_pat_cur_offset_2 + _source_stream_max_pool_serial_6_source_1_pat_cur_offset_3;
  wire _set_flag_1209;
  assign _set_flag_1209 = max_pool_serial_6_comp_fsm == 4;
  reg _tmp_1210;
  reg _tmp_1211;
  reg _tmp_1212;
  reg _tmp_1213;
  reg _tmp_1214;
  reg _tmp_1215;
  reg _tmp_1216;
  localparam _tmp_1217 = 33;
  wire [_tmp_1217-1:0] _tmp_1218;
  assign _tmp_1218 = max_pool_serial_6_stream_out_local + max_pool_serial_6_out_page_comp_offset_buf;
  reg [_tmp_1217-1:0] _tmp_1219;
  reg [_tmp_1217-1:0] _tmp_1220;
  reg [_tmp_1217-1:0] _tmp_1221;
  reg [_tmp_1217-1:0] _tmp_1222;
  reg [_tmp_1217-1:0] _tmp_1223;
  reg [_tmp_1217-1:0] _tmp_1224;
  reg [_tmp_1217-1:0] _tmp_1225;
  reg [6-1:0] _tmp_1226;
  reg [6-1:0] _tmp_1227;
  reg [6-1:0] _tmp_1228;
  reg [6-1:0] _tmp_1229;
  reg [6-1:0] _tmp_1230;
  reg [6-1:0] _tmp_1231;
  reg [6-1:0] _tmp_1232;
  wire [1-1:0] write_rtl_bank_1233;
  assign write_rtl_bank_1233 = _stream_max_pool_serial_6_sink_5_sink_waddr;
  assign ram_w16_l8192_id0_0_0_wdata = (_stream_max_pool_serial_6_stream_oready && _stream_max_pool_serial_6_sink_5_sink_wenable && (_stream_max_pool_serial_6_sink_5_sink_sel == 2) && (write_rtl_bank_1233 == 0))? _stream_max_pool_serial_6_sink_5_sink_wdata : 'hx;
  assign ram_w16_l8192_id0_0_0_wenable = (_stream_max_pool_serial_6_stream_oready && _stream_max_pool_serial_6_sink_5_sink_wenable && (_stream_max_pool_serial_6_sink_5_sink_sel == 2) && (write_rtl_bank_1233 == 0))? 1'd1 : 0;
  assign ram_w16_l8192_id0_1_0_wdata = (_stream_max_pool_serial_6_stream_oready && _stream_max_pool_serial_6_sink_5_sink_wenable && (_stream_max_pool_serial_6_sink_5_sink_sel == 2) && (write_rtl_bank_1233 == 1))? _stream_max_pool_serial_6_sink_5_sink_wdata : 'hx;
  assign ram_w16_l8192_id0_1_0_wenable = (_stream_max_pool_serial_6_stream_oready && _stream_max_pool_serial_6_sink_5_sink_wenable && (_stream_max_pool_serial_6_sink_5_sink_sel == 2) && (write_rtl_bank_1233 == 1))? 1'd1 : 0;
  reg [32-1:0] _stream_max_pool_serial_6_sink_5_sink_fsm_1;
  localparam _stream_max_pool_serial_6_sink_5_sink_fsm_1_init = 0;
  wire _set_flag_1234;
  assign _set_flag_1234 = max_pool_serial_6_comp_fsm == 5;
  assign _stream_max_pool_serial_6_run_flag = (_set_flag_1234)? 1 : 0;
  reg _tmp_1235;
  reg _tmp_1236;
  reg _tmp_1237;
  reg _tmp_1238;
  reg _tmp_1239;
  reg _tmp_1240;
  reg _tmp_1241;
  reg _tmp_1242;
  reg _tmp_1243;
  reg _tmp_1244;
  assign __reduce_max_27_source_stop = __reduce_max_27_stream_oready && 1'd0;
  reg _tmp_1245;
  reg _tmp_1246;
  reg _tmp_1247;
  assign __reduce_max_27_sink_start = _tmp_1247;
  reg _tmp_1248;
  reg _tmp_1249;
  reg _tmp_1250;
  assign __reduce_max_27_sink_stop = _tmp_1250;
  reg _tmp_1251;
  reg _tmp_1252;
  reg _tmp_1253;
  assign __reduce_max_27_sink_busy = _tmp_1253;
  reg _tmp_1254;
  assign __reduce_max_27_busy = __reduce_max_27_source_busy || __reduce_max_27_sink_busy || __reduce_max_27_busy_reg;
  reg _tmp_1255;
  reg _tmp_1256;
  reg _tmp_1257;
  reg _tmp_1258;
  reg _tmp_1259;
  reg _tmp_1260;
  reg [1-1:0] __variable_wdata_2140;
  assign stream_max_pool_serial_6__reduce_reset_data = __variable_wdata_2140;
  reg _tmp_1261;
  reg _tmp_1262;
  reg _tmp_1263;
  reg _tmp_1264;
  assign _stream_max_pool_serial_6_source_stop = _stream_max_pool_serial_6_stream_oready && (_stream_max_pool_serial_6_source_1_idle && (_stream_max_pool_serial_6_fsm == 3));
  localparam _tmp_1265 = 1;
  wire [_tmp_1265-1:0] _tmp_1266;
  assign _tmp_1266 = _stream_max_pool_serial_6_source_1_idle && (_stream_max_pool_serial_6_fsm == 3);
  reg [_tmp_1265-1:0] _tmp_1267;
  localparam _tmp_1268 = 1;
  wire [_tmp_1268-1:0] _tmp_1269;
  assign _tmp_1269 = _stream_max_pool_serial_6_source_1_idle && (_stream_max_pool_serial_6_fsm == 3);
  reg [_tmp_1268-1:0] _tmp_1270;
  reg _tmp_1271;
  reg _tmp_1272;
  reg _tmp_1273;
  reg _tmp_1274;
  reg _tmp_1275;
  reg _tmp_1276;
  reg _tmp_1277;
  assign _stream_max_pool_serial_6_sink_start = _tmp_1277;
  reg _tmp_1278;
  reg _tmp_1279;
  reg _tmp_1280;
  reg _tmp_1281;
  reg _tmp_1282;
  reg _tmp_1283;
  reg _tmp_1284;
  assign _stream_max_pool_serial_6_sink_stop = _tmp_1284;
  reg _tmp_1285;
  reg _tmp_1286;
  reg _tmp_1287;
  reg _tmp_1288;
  reg _tmp_1289;
  reg _tmp_1290;
  reg _tmp_1291;
  assign _stream_max_pool_serial_6_sink_busy = _tmp_1291;
  reg _tmp_1292;
  assign _stream_max_pool_serial_6_busy = _stream_max_pool_serial_6_source_busy || _stream_max_pool_serial_6_sink_busy || _stream_max_pool_serial_6_busy_reg;
  wire [9-1:0] _dma_write_packed_high_local_size_1293;
  assign _dma_write_packed_high_local_size_1293 = cparam_max_pool_serial_6_out_write_size >> 1;
  wire [1-1:0] _dma_write_packed_low_local_size_1294;
  assign _dma_write_packed_low_local_size_1294 = cparam_max_pool_serial_6_out_write_size & { 1{ 1'd1 } };
  wire [9-1:0] _dma_write_packed_local_packed_size_1295;
  assign _dma_write_packed_local_packed_size_1295 = (_dma_write_packed_low_local_size_1294 > 0)? _dma_write_packed_high_local_size_1293 + 1 : _dma_write_packed_high_local_size_1293;
  wire [32-1:0] mask_addr_shifted_1296;
  assign mask_addr_shifted_1296 = max_pool_serial_6_objaddr + max_pool_serial_6_out_base_offset + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_1297;
  assign mask_addr_masked_1297 = mask_addr_shifted_1296 << 2;
  reg [32-1:0] read_burst_packed_fsm_57;
  localparam read_burst_packed_fsm_57_init = 0;
  reg [13-1:0] read_burst_packed_addr_1298;
  reg [13-1:0] read_burst_packed_stride_1299;
  reg [33-1:0] read_burst_packed_length_1300;
  reg read_burst_packed_rvalid_1301;
  reg read_burst_packed_rlast_1302;
  wire [12-1:0] read_burst_packed_ram_addr_1303;
  assign read_burst_packed_ram_addr_1303 = read_burst_packed_addr_1298 >> 1;
  localparam _tmp_1304 = 1;
  wire [_tmp_1304-1:0] _tmp_1305;
  assign _tmp_1305 = (read_burst_packed_fsm_57 == 1) && (!read_burst_packed_rvalid_1301 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0));
  reg [_tmp_1304-1:0] __tmp_1305_1;
  wire [16-1:0] read_burst_packed_ram_rdata_1306;
  assign read_burst_packed_ram_rdata_1306 = ram_w16_l8192_id0_0_1_rdata;
  wire [12-1:0] read_burst_packed_ram_addr_1307;
  assign read_burst_packed_ram_addr_1307 = read_burst_packed_addr_1298 >> 1;
  localparam _tmp_1308 = 1;
  wire [_tmp_1308-1:0] _tmp_1309;
  assign _tmp_1309 = (read_burst_packed_fsm_57 == 1) && (!read_burst_packed_rvalid_1301 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0));
  reg [_tmp_1308-1:0] __tmp_1309_1;
  wire [16-1:0] read_burst_packed_ram_rdata_1310;
  assign read_burst_packed_ram_rdata_1310 = ram_w16_l8192_id0_1_1_rdata;
  wire [32-1:0] read_burst_packed_rdata_1311;
  assign read_burst_packed_rdata_1311 = { read_burst_packed_ram_rdata_1310, read_burst_packed_ram_rdata_1306 };
  reg _maxi_wdata_cond_1_1;
  reg [32-1:0] matmul_11_objaddr;
  reg [32-1:0] matmul_11_arg_objaddr_0;
  reg [32-1:0] matmul_11_arg_objaddr_1;
  reg [32-1:0] matmul_11_arg_objaddr_2;
  reg [32-1:0] matmul_11_arg_objaddr_3;
  reg [32-1:0] control_matmul_11;
  localparam control_matmul_11_init = 0;
  reg _control_matmul_11_called;
  wire signed [32-1:0] matmul_11_act_base_offset;
  reg signed [32-1:0] matmul_11_act_base_offset_row;
  reg signed [32-1:0] matmul_11_act_base_offset_bat;
  assign matmul_11_act_base_offset = matmul_11_act_base_offset_row + matmul_11_act_base_offset_bat;
  reg signed [32-1:0] matmul_11_filter_base_offset;
  reg [32-1:0] matmul_11_next_stream_num_ops;
  wire signed [32-1:0] matmul_11_out_base_offset;
  reg signed [32-1:0] matmul_11_out_base_offset_val;
  reg signed [32-1:0] matmul_11_out_base_offset_col;
  reg signed [32-1:0] matmul_11_out_base_offset_row;
  reg signed [32-1:0] matmul_11_out_base_offset_bat;
  reg signed [32-1:0] matmul_11_out_base_offset_och;
  assign matmul_11_out_base_offset = matmul_11_out_base_offset_val + matmul_11_out_base_offset_col + matmul_11_out_base_offset_row + matmul_11_out_base_offset_bat + matmul_11_out_base_offset_och;
  reg matmul_11_dma_flag_0;
  reg [32-1:0] matmul_11_sync_comp_count;
  reg [32-1:0] matmul_11_sync_out_count;
  reg [32-1:0] matmul_11_write_count;
  reg [32-1:0] matmul_11_next_out_write_size;
  reg [32-1:0] matmul_11_col_count;
  reg [32-1:0] matmul_11_row_count;
  reg [32-1:0] matmul_11_bat_count;
  reg [32-1:0] matmul_11_och_count;
  reg [1-1:0] matmul_11_col_select;
  reg [1-1:0] matmul_11_row_select;
  reg [32-1:0] matmul_11_out_col_count;
  reg [32-1:0] matmul_11_out_row_count;
  reg [32-1:0] matmul_11_out_ram_select;
  reg [32-1:0] matmul_11_prev_col_count;
  reg [32-1:0] matmul_11_prev_row_count;
  reg [32-1:0] matmul_11_prev_bat_count;
  reg [32-1:0] matmul_11_prev_och_count;
  reg [1-1:0] matmul_11_prev_row_select;
  reg [32-1:0] matmul_11_stream_act_local_0;
  reg [32-1:0] matmul_11_stream_out_local_val;
  reg [32-1:0] matmul_11_stream_out_local_col;
  wire [32-1:0] matmul_11_stream_out_local;
  assign matmul_11_stream_out_local = matmul_11_stream_out_local_val + matmul_11_stream_out_local_col;
  reg [32-1:0] matmul_11_act_page_comp_offset_0;
  reg [32-1:0] matmul_11_act_page_dma_offset_0;
  reg [32-1:0] matmul_11_filter_page_comp_offset;
  reg [32-1:0] matmul_11_filter_page_dma_offset;
  reg matmul_11_out_page;
  reg [32-1:0] matmul_11_out_page_comp_offset;
  reg [32-1:0] matmul_11_out_page_dma_offset;
  reg [32-1:0] matmul_11_out_laddr_offset;
  reg matmul_11_skip_read_filter;
  reg matmul_11_skip_read_act;
  reg matmul_11_skip_comp;
  reg matmul_11_skip_write_out;
  wire [8-1:0] _dma_read_packed_high_local_size_1312;
  assign _dma_read_packed_high_local_size_1312 = cparam_matmul_11_bias_num >> 1;
  wire [1-1:0] _dma_read_packed_low_local_size_1313;
  assign _dma_read_packed_low_local_size_1313 = cparam_matmul_11_bias_num & { 1{ 1'd1 } };
  wire [8-1:0] _dma_read_packed_local_packed_size_1314;
  assign _dma_read_packed_local_packed_size_1314 = (_dma_read_packed_low_local_size_1313 > 0)? _dma_read_packed_high_local_size_1312 + 1 : _dma_read_packed_high_local_size_1312;
  wire [32-1:0] mask_addr_shifted_1315;
  assign mask_addr_shifted_1315 = matmul_11_arg_objaddr_2 + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_1316;
  assign mask_addr_masked_1316 = mask_addr_shifted_1315 << 2;
  reg [32-1:0] write_burst_packed_fsm_58;
  localparam write_burst_packed_fsm_58_init = 0;
  reg [9-1:0] write_burst_packed_addr_1317;
  reg [9-1:0] write_burst_packed_stride_1318;
  reg [33-1:0] write_burst_packed_length_1319;
  reg write_burst_packed_done_1320;
  wire [8-1:0] write_burst_packed_ram_addr_1321;
  assign write_burst_packed_ram_addr_1321 = write_burst_packed_addr_1317 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_1322;
  assign write_burst_packed_ram_wdata_1322 = _maxi_rdata_sb_0 >> 0;
  assign ram_w16_l512_id1_0_1_addr = ((write_burst_packed_fsm_58 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_addr_1321 : 
                                     ((write_burst_packed_fsm_34 == 1) && write_burst_block_ram_wvalid_118)? write_burst_packed_ram_addr_124 : 'hx;
  assign ram_w16_l512_id1_0_1_wdata = ((write_burst_packed_fsm_58 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_wdata_1322 : 
                                      ((write_burst_packed_fsm_34 == 1) && write_burst_block_ram_wvalid_118)? write_burst_packed_ram_wdata_125 : 'hx;
  assign ram_w16_l512_id1_0_1_wenable = ((write_burst_packed_fsm_58 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 
                                        ((write_burst_packed_fsm_34 == 1) && write_burst_block_ram_wvalid_118)? 1'd1 : 0;
  assign ram_w16_l512_id1_0_1_enable = ((write_burst_packed_fsm_58 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 
                                       ((write_burst_packed_fsm_34 == 1) && write_burst_block_ram_wvalid_118)? 1'd1 : 0;
  wire [8-1:0] write_burst_packed_ram_addr_1323;
  assign write_burst_packed_ram_addr_1323 = write_burst_packed_addr_1317 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_1324;
  assign write_burst_packed_ram_wdata_1324 = _maxi_rdata_sb_0 >> 16;
  assign ram_w16_l512_id1_1_1_addr = ((write_burst_packed_fsm_58 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_addr_1323 : 
                                     ((write_burst_packed_fsm_34 == 1) && write_burst_block_ram_wvalid_118)? write_burst_packed_ram_addr_126 : 'hx;
  assign ram_w16_l512_id1_1_1_wdata = ((write_burst_packed_fsm_58 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_wdata_1324 : 
                                      ((write_burst_packed_fsm_34 == 1) && write_burst_block_ram_wvalid_118)? write_burst_packed_ram_wdata_127 : 'hx;
  assign ram_w16_l512_id1_1_1_wenable = ((write_burst_packed_fsm_58 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 
                                        ((write_burst_packed_fsm_34 == 1) && write_burst_block_ram_wvalid_118)? 1'd1 : 0;
  assign ram_w16_l512_id1_1_1_enable = ((write_burst_packed_fsm_58 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 
                                       ((write_burst_packed_fsm_34 == 1) && write_burst_block_ram_wvalid_118)? 1'd1 : 0;
  wire [8-1:0] _dma_read_packed_high_local_size_1325;
  assign _dma_read_packed_high_local_size_1325 = cparam_matmul_11_scale_num >> 1;
  wire [1-1:0] _dma_read_packed_low_local_size_1326;
  assign _dma_read_packed_low_local_size_1326 = cparam_matmul_11_scale_num & { 1{ 1'd1 } };
  wire [8-1:0] _dma_read_packed_local_packed_size_1327;
  assign _dma_read_packed_local_packed_size_1327 = (_dma_read_packed_low_local_size_1326 > 0)? _dma_read_packed_high_local_size_1325 + 1 : _dma_read_packed_high_local_size_1325;
  wire [32-1:0] mask_addr_shifted_1328;
  assign mask_addr_shifted_1328 = matmul_11_arg_objaddr_3 + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_1329;
  assign mask_addr_masked_1329 = mask_addr_shifted_1328 << 2;
  reg [32-1:0] write_burst_packed_fsm_59;
  localparam write_burst_packed_fsm_59_init = 0;
  reg [9-1:0] write_burst_packed_addr_1330;
  reg [9-1:0] write_burst_packed_stride_1331;
  reg [33-1:0] write_burst_packed_length_1332;
  reg write_burst_packed_done_1333;
  wire [8-1:0] write_burst_packed_ram_addr_1334;
  assign write_burst_packed_ram_addr_1334 = write_burst_packed_addr_1330 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_1335;
  assign write_burst_packed_ram_wdata_1335 = _maxi_rdata_sb_0 >> 0;
  assign ram_w16_l512_id2_0_1_addr = ((write_burst_packed_fsm_59 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_addr_1334 : 
                                     ((write_burst_packed_fsm_35 == 1) && write_burst_block_ram_wvalid_128)? write_burst_packed_ram_addr_134 : 'hx;
  assign ram_w16_l512_id2_0_1_wdata = ((write_burst_packed_fsm_59 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_wdata_1335 : 
                                      ((write_burst_packed_fsm_35 == 1) && write_burst_block_ram_wvalid_128)? write_burst_packed_ram_wdata_135 : 'hx;
  assign ram_w16_l512_id2_0_1_wenable = ((write_burst_packed_fsm_59 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 
                                        ((write_burst_packed_fsm_35 == 1) && write_burst_block_ram_wvalid_128)? 1'd1 : 0;
  assign ram_w16_l512_id2_0_1_enable = ((write_burst_packed_fsm_59 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 
                                       ((write_burst_packed_fsm_35 == 1) && write_burst_block_ram_wvalid_128)? 1'd1 : 0;
  wire [8-1:0] write_burst_packed_ram_addr_1336;
  assign write_burst_packed_ram_addr_1336 = write_burst_packed_addr_1330 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_1337;
  assign write_burst_packed_ram_wdata_1337 = _maxi_rdata_sb_0 >> 16;
  assign ram_w16_l512_id2_1_1_addr = ((write_burst_packed_fsm_59 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_addr_1336 : 
                                     ((write_burst_packed_fsm_35 == 1) && write_burst_block_ram_wvalid_128)? write_burst_packed_ram_addr_136 : 'hx;
  assign ram_w16_l512_id2_1_1_wdata = ((write_burst_packed_fsm_59 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_wdata_1337 : 
                                      ((write_burst_packed_fsm_35 == 1) && write_burst_block_ram_wvalid_128)? write_burst_packed_ram_wdata_137 : 'hx;
  assign ram_w16_l512_id2_1_1_wenable = ((write_burst_packed_fsm_59 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 
                                        ((write_burst_packed_fsm_35 == 1) && write_burst_block_ram_wvalid_128)? 1'd1 : 0;
  assign ram_w16_l512_id2_1_1_enable = ((write_burst_packed_fsm_59 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 
                                       ((write_burst_packed_fsm_35 == 1) && write_burst_block_ram_wvalid_128)? 1'd1 : 0;
  wire [14-1:0] _dma_read_packed_high_local_size_1338;
  assign _dma_read_packed_high_local_size_1338 = cparam_matmul_11_filter_read_size >> 1;
  wire [1-1:0] _dma_read_packed_low_local_size_1339;
  assign _dma_read_packed_low_local_size_1339 = cparam_matmul_11_filter_read_size & { 1{ 1'd1 } };
  wire [14-1:0] _dma_read_packed_local_packed_size_1340;
  assign _dma_read_packed_local_packed_size_1340 = (_dma_read_packed_low_local_size_1339 > 0)? _dma_read_packed_high_local_size_1338 + 1 : _dma_read_packed_high_local_size_1338;
  wire [32-1:0] mask_addr_shifted_1341;
  assign mask_addr_shifted_1341 = matmul_11_arg_objaddr_1 + matmul_11_filter_base_offset + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_1342;
  assign mask_addr_masked_1342 = mask_addr_shifted_1341 << 2;
  wire [32-1:0] matmul_11_mux_act_gaddr_0;
  assign matmul_11_mux_act_gaddr_0 = (matmul_11_row_select == 0)? matmul_11_arg_objaddr_0 + (matmul_11_act_base_offset + cparam_matmul_11_act_offset_values_0) : 1'd0;
  wire matmul_11_dma_pad_mask_0;
  assign matmul_11_dma_pad_mask_0 = (matmul_11_row_count + 0 < cparam_matmul_11_pad_row_top) || (matmul_11_row_count + 0 >= cparam_matmul_11_act_num_row + cparam_matmul_11_pad_row_top);
  wire matmul_11_mux_dma_pad_mask_0;
  assign matmul_11_mux_dma_pad_mask_0 = (matmul_11_row_select == 0)? matmul_11_dma_pad_mask_0 : 1'd0;
  wire matmul_11_mux_dma_flag_0;
  assign matmul_11_mux_dma_flag_0 = (matmul_11_prev_row_select == 0)? matmul_11_dma_flag_0 : 1'd0;
  wire [13-1:0] _dma_read_packed_high_local_size_1343;
  assign _dma_read_packed_high_local_size_1343 = cparam_matmul_11_act_read_size >> 1;
  wire [1-1:0] _dma_read_packed_low_local_size_1344;
  assign _dma_read_packed_low_local_size_1344 = cparam_matmul_11_act_read_size & { 1{ 1'd1 } };
  wire [13-1:0] _dma_read_packed_local_packed_size_1345;
  assign _dma_read_packed_local_packed_size_1345 = (_dma_read_packed_low_local_size_1344 > 0)? _dma_read_packed_high_local_size_1343 + 1 : _dma_read_packed_high_local_size_1343;
  wire [32-1:0] mask_addr_shifted_1346;
  assign mask_addr_shifted_1346 = matmul_11_mux_act_gaddr_0 + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_1347;
  assign mask_addr_masked_1347 = mask_addr_shifted_1346 << 2;
  assign _maxi_read_req_fifo_deq = ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 10)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 9)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 8)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 7)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 6)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 5)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 4)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 3)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 2)) && !_maxi_read_req_fifo_empty)? 1 : 
                                   ((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 1)) && !_maxi_read_req_fifo_empty)? 1 : 0;
  reg [32-1:0] write_burst_packed_fsm_60;
  localparam write_burst_packed_fsm_60_init = 0;
  reg [13-1:0] write_burst_packed_addr_1348;
  reg [13-1:0] write_burst_packed_stride_1349;
  reg [33-1:0] write_burst_packed_length_1350;
  reg write_burst_packed_done_1351;
  wire [12-1:0] write_burst_packed_ram_addr_1352;
  assign write_burst_packed_ram_addr_1352 = write_burst_packed_addr_1348 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_1353;
  assign write_burst_packed_ram_wdata_1353 = _maxi_rdata_sb_0 >> 0;
  assign ram_w16_l8192_id0_0_1_addr = ((write_burst_packed_fsm_60 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_addr_1352 : 
                                      ((read_burst_packed_fsm_57 == 1) && (!read_burst_packed_rvalid_1301 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? read_burst_packed_ram_addr_1303 : 'hx;
  assign ram_w16_l8192_id0_0_1_wdata = ((write_burst_packed_fsm_60 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_wdata_1353 : 'hx;
  assign ram_w16_l8192_id0_0_1_wenable = ((write_burst_packed_fsm_60 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  assign ram_w16_l8192_id0_0_1_enable = ((write_burst_packed_fsm_60 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 
                                        ((read_burst_packed_fsm_57 == 1) && (!read_burst_packed_rvalid_1301 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? 1'd1 : 0;
  wire [12-1:0] write_burst_packed_ram_addr_1354;
  assign write_burst_packed_ram_addr_1354 = write_burst_packed_addr_1348 >> 1;
  wire [16-1:0] write_burst_packed_ram_wdata_1355;
  assign write_burst_packed_ram_wdata_1355 = _maxi_rdata_sb_0 >> 16;
  assign ram_w16_l8192_id0_1_1_addr = ((write_burst_packed_fsm_60 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_addr_1354 : 
                                      ((read_burst_packed_fsm_57 == 1) && (!read_burst_packed_rvalid_1301 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? read_burst_packed_ram_addr_1307 : 'hx;
  assign ram_w16_l8192_id0_1_1_wdata = ((write_burst_packed_fsm_60 == 1) && _maxi_rvalid_sb_0)? write_burst_packed_ram_wdata_1355 : 'hx;
  assign ram_w16_l8192_id0_1_1_wenable = ((write_burst_packed_fsm_60 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 0;
  assign ram_w16_l8192_id0_1_1_enable = ((write_burst_packed_fsm_60 == 1) && _maxi_rvalid_sb_0)? 1'd1 : 
                                        ((read_burst_packed_fsm_57 == 1) && (!read_burst_packed_rvalid_1301 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? 1'd1 : 0;
  assign _maxi_rready_sb_0 = (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2) || (_maxi_read_data_fsm == 2);
  reg [32-1:0] matmul_11_comp_fsm;
  localparam matmul_11_comp_fsm_init = 0;
  reg [32-1:0] matmul_11_filter_page_comp_offset_buf;
  reg [32-1:0] matmul_11_act_page_comp_offset_buf_0;
  reg [32-1:0] matmul_11_out_page_comp_offset_buf;
  reg [32-1:0] matmul_11_row_count_buf;
  reg [1-1:0] matmul_11_row_select_buf;
  reg [32-1:0] matmul_11_och_count_buf;
  wire matmul_11_stream_pad_mask_0_0;
  assign matmul_11_stream_pad_mask_0_0 = (matmul_11_col_count + 0 < cparam_matmul_11_pad_col_left) || (matmul_11_col_count + 0 >= cparam_matmul_11_act_num_col + cparam_matmul_11_pad_col_left) || (matmul_11_row_count_buf + 0 < cparam_matmul_11_pad_row_top) || (matmul_11_row_count_buf + 0 >= cparam_matmul_11_act_num_row + cparam_matmul_11_pad_row_top);
  reg [1-1:0] matmul_11_stream_pad_masks;
  wire [13-1:0] stream_matmul_11_parameter_0_data;
  wire [1-1:0] stream_matmul_11_parameter_1_data;
  wire [1-1:0] stream_matmul_11_parameter_2_data;
  wire [1-1:0] stream_matmul_11_parameter_3_data;
  wire [1-1:0] stream_matmul_11_parameter_4_data;
  wire [1-1:0] stream_matmul_11__reduce_reset_data;
  wire [1-1:0] stream_matmul_11_parameter_6_data;
  wire [16-1:0] stream_matmul_11_source_7_data;
  wire [1-1:0] stream_matmul_11_parameter_8_data;
  wire [16-1:0] stream_matmul_11_source_9_data;
  wire [1-1:0] stream_matmul_11_parameter_10_data;
  wire [16-1:0] stream_matmul_11_source_11_data;
  wire [1-1:0] stream_matmul_11_parameter_12_data;
  wire [16-1:0] stream_matmul_11_source_13_data;
  wire [1-1:0] stream_matmul_11_parameter_14_data;
  wire [16-1:0] stream_matmul_11_source_15_data;
  wire [1-1:0] stream_matmul_11_parameter_16_data;
  wire [1-1:0] stream_matmul_11_parameter_17_data;
  wire [5-1:0] stream_matmul_11_parameter_18_data;
  wire [2-1:0] stream_matmul_11_parameter_19_data;
  wire [16-1:0] stream_matmul_11_source_20_data;
  wire [16-1:0] stream_matmul_11_source_21_data;
  reg __stream_matmul_11_stream_ivalid_1;
  reg __stream_matmul_11_stream_ivalid_2;
  reg __stream_matmul_11_stream_ivalid_3;
  reg __stream_matmul_11_stream_ivalid_4;
  reg __stream_matmul_11_stream_ivalid_5;
  reg __stream_matmul_11_stream_ivalid_6;
  reg __stream_matmul_11_stream_ivalid_7;
  reg __stream_matmul_11_stream_ivalid_8;
  reg __stream_matmul_11_stream_ivalid_9;
  reg __stream_matmul_11_stream_ivalid_10;
  reg __stream_matmul_11_stream_ivalid_11;
  reg __stream_matmul_11_stream_ivalid_12;
  reg __stream_matmul_11_stream_ivalid_13;
  reg __stream_matmul_11_stream_ivalid_14;
  reg __stream_matmul_11_stream_ivalid_15;
  reg __stream_matmul_11_stream_ivalid_16;
  reg __stream_matmul_11_stream_ivalid_17;
  reg __stream_matmul_11_stream_ivalid_18;
  reg __stream_matmul_11_stream_ivalid_19;
  reg __stream_matmul_11_stream_ivalid_20;
  reg __stream_matmul_11_stream_ivalid_21;
  reg __stream_matmul_11_stream_ivalid_22;
  reg __stream_matmul_11_stream_ivalid_23;
  reg __stream_matmul_11_stream_ivalid_24;
  reg __stream_matmul_11_stream_ivalid_25;
  reg __stream_matmul_11_stream_ivalid_26;
  reg __stream_matmul_11_stream_ivalid_27;
  reg __stream_matmul_11_stream_ivalid_28;
  reg __stream_matmul_11_stream_ivalid_29;
  wire [16-1:0] _slice_data_2175;
  assign _slice_data_2175 = stream_matmul_11_source_7_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_2176;
  assign _reinterpretcast_src_2176 = _slice_data_2175;
  wire signed [16-1:0] _reinterpretcast_data_2176;
  assign _reinterpretcast_data_2176 = _reinterpretcast_src_2176;
  wire signed [16-1:0] _cond_data_2177;
  assign _cond_data_2177 = (stream_matmul_11_parameter_6_data)? _reinterpretcast_data_2176 : _reinterpretcast_data_2176;
  wire [16-1:0] _slice_data_2182;
  assign _slice_data_2182 = stream_matmul_11_source_9_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_2183;
  assign _reinterpretcast_src_2183 = _slice_data_2182;
  wire signed [16-1:0] _reinterpretcast_data_2183;
  assign _reinterpretcast_data_2183 = _reinterpretcast_src_2183;
  wire signed [16-1:0] _cond_data_2184;
  assign _cond_data_2184 = (stream_matmul_11_parameter_8_data)? _reinterpretcast_data_2183 : _reinterpretcast_data_2183;
  wire [16-1:0] _slice_data_2189;
  assign _slice_data_2189 = stream_matmul_11_source_11_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_2190;
  assign _reinterpretcast_src_2190 = _slice_data_2189;
  wire [16-1:0] _reinterpretcast_data_2190;
  assign _reinterpretcast_data_2190 = _reinterpretcast_src_2190;
  wire [16-1:0] _cond_data_2191;
  assign _cond_data_2191 = (stream_matmul_11_parameter_10_data)? _reinterpretcast_data_2190 : _reinterpretcast_data_2190;
  wire [16-1:0] _slice_data_2196;
  assign _slice_data_2196 = stream_matmul_11_source_13_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_2197;
  assign _reinterpretcast_src_2197 = _slice_data_2196;
  wire [16-1:0] _reinterpretcast_data_2197;
  assign _reinterpretcast_data_2197 = _reinterpretcast_src_2197;
  wire [16-1:0] _cond_data_2198;
  assign _cond_data_2198 = (stream_matmul_11_parameter_12_data)? _reinterpretcast_data_2197 : _reinterpretcast_data_2197;
  wire [16-1:0] _slice_data_2203;
  assign _slice_data_2203 = stream_matmul_11_source_15_data[5'd15:1'd0];
  wire [16-1:0] _reinterpretcast_src_2204;
  assign _reinterpretcast_src_2204 = _slice_data_2203;
  wire [16-1:0] _reinterpretcast_data_2204;
  assign _reinterpretcast_data_2204 = _reinterpretcast_src_2204;
  wire [16-1:0] _cond_data_2205;
  assign _cond_data_2205 = (stream_matmul_11_parameter_14_data)? _reinterpretcast_data_2204 : _reinterpretcast_data_2204;
  reg [1-1:0] _eq_data_2211;
  reg [1-1:0] _eq_data_2215;
  wire [16-1:0] _reinterpretcast_src_2229;
  assign _reinterpretcast_src_2229 = stream_matmul_11_source_21_data;
  wire signed [16-1:0] _reinterpretcast_data_2229;
  assign _reinterpretcast_data_2229 = _reinterpretcast_src_2229;
  wire [1-1:0] _pointer_data_2230;
  assign _pointer_data_2230 = stream_matmul_11_parameter_3_data[1'sd0];
  reg [16-1:0] _plus_data_2235;
  reg [16-1:0] _plus_data_2240;
  reg [16-1:0] _plus_data_2245;
  reg [1-1:0] _eq_data_2251;
  reg [1-1:0] _eq_data_2254;
  reg [16-1:0] __delay_data_2403__variable_2210;
  reg [1-1:0] __delay_data_2404_pointer_2230;
  reg signed [16-1:0] __delay_data_2405_reinterpretcast_2229;
  reg [1-1:0] __delay_data_2406__variable_2161;
  reg [13-1:0] __delay_data_2427__variable_2156;
  reg signed [16-1:0] __delay_data_2438_cond_2177;
  reg signed [16-1:0] __delay_data_2455_cond_2184;
  wire signed [16-1:0] _cond_data_2213;
  assign _cond_data_2213 = (_eq_data_2211)? __delay_data_2403__variable_2210 : 1'sd0;
  wire signed [16-1:0] _cond_data_2217;
  assign _cond_data_2217 = (_eq_data_2215)? _cond_data_2213 : 1'sd0;
  wire signed [16-1:0] _reinterpretcast_src_2223;
  assign _reinterpretcast_src_2223 = _cond_data_2217;
  wire signed [16-1:0] _reinterpretcast_data_2223;
  assign _reinterpretcast_data_2223 = _reinterpretcast_src_2223;
  wire signed [16-1:0] _cond_data_2233;
  assign _cond_data_2233 = (__delay_data_2404_pointer_2230)? 1'sd0 : _reinterpretcast_data_2223;
  assign _mul_18_is_root = ((_stream_matmul_11_busy)? 0 : 1) && (((_stream_conv2d_4_busy)? 0 : 1) && 1);
  assign _mul_18_stream_oready = ((_stream_matmul_11_busy)? _stream_matmul_11_stream_oready : 1) && (((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_18_stream_internal_oready);
  reg [1-1:0] __delay_data_2407__delay_2406__variable_2161;
  reg [16-1:0] __delay_data_2417_plus_2240;
  reg [13-1:0] __delay_data_2428__delay_2427__variable_2156;
  reg signed [16-1:0] __delay_data_2439__delay_2438_cond_2177;
  reg signed [16-1:0] __delay_data_2456__delay_2455_cond_2184;
  reg [16-1:0] __delay_data_2473_plus_2245;
  reg [1-1:0] __delay_data_2491_eq_2251;
  reg [1-1:0] __delay_data_2520_eq_2254;
  reg [1-1:0] __delay_data_2408__delay_2407__delay_2406__variable_2161;
  reg [16-1:0] __delay_data_2418__delay_2417_plus_2240;
  reg [13-1:0] __delay_data_2429__delay_2428__delay_2427__variable_2156;
  reg signed [16-1:0] __delay_data_2440__delay_2439__delay_2438_cond_2177;
  reg signed [16-1:0] __delay_data_2457__delay_2456__delay_2455_cond_2184;
  reg [16-1:0] __delay_data_2474__delay_2473_plus_2245;
  reg [1-1:0] __delay_data_2492__delay_2491_eq_2251;
  reg [1-1:0] __delay_data_2521__delay_2520_eq_2254;
  reg [1-1:0] __delay_data_2409__delay_2408__delay_2407____variable_2161;
  reg [16-1:0] __delay_data_2419__delay_2418__delay_2417_plus_2240;
  reg [13-1:0] __delay_data_2430__delay_2429__delay_2428____variable_2156;
  reg signed [16-1:0] __delay_data_2441__delay_2440__delay_2439___cond_2177;
  reg signed [16-1:0] __delay_data_2458__delay_2457__delay_2456___cond_2184;
  reg [16-1:0] __delay_data_2475__delay_2474__delay_2473_plus_2245;
  reg [1-1:0] __delay_data_2493__delay_2492__delay_2491_eq_2251;
  reg [1-1:0] __delay_data_2522__delay_2521__delay_2520_eq_2254;
  reg [1-1:0] __delay_data_2410__delay_2409__delay_2408____variable_2161;
  reg [16-1:0] __delay_data_2420__delay_2419__delay_2418___plus_2240;
  reg [13-1:0] __delay_data_2431__delay_2430__delay_2429____variable_2156;
  reg signed [16-1:0] __delay_data_2442__delay_2441__delay_2440___cond_2177;
  reg signed [16-1:0] __delay_data_2459__delay_2458__delay_2457___cond_2184;
  reg [16-1:0] __delay_data_2476__delay_2475__delay_2474___plus_2245;
  reg [1-1:0] __delay_data_2494__delay_2493__delay_2492__delay_2491_eq_2251;
  reg [1-1:0] __delay_data_2523__delay_2522__delay_2521__delay_2520_eq_2254;
  reg [1-1:0] __delay_data_2411__delay_2410__delay_2409____variable_2161;
  reg [16-1:0] __delay_data_2421__delay_2420__delay_2419___plus_2240;
  reg [13-1:0] __delay_data_2432__delay_2431__delay_2430____variable_2156;
  reg signed [16-1:0] __delay_data_2443__delay_2442__delay_2441___cond_2177;
  reg signed [16-1:0] __delay_data_2460__delay_2459__delay_2458___cond_2184;
  reg [16-1:0] __delay_data_2477__delay_2476__delay_2475___plus_2245;
  reg [1-1:0] __delay_data_2495__delay_2494__delay_2493__delay_2492___eq_2251;
  reg [1-1:0] __delay_data_2524__delay_2523__delay_2522__delay_2521___eq_2254;
  reg [1-1:0] __delay_data_2412__delay_2411__delay_2410____variable_2161;
  reg [16-1:0] __delay_data_2422__delay_2421__delay_2420___plus_2240;
  reg [13-1:0] __delay_data_2433__delay_2432__delay_2431____variable_2156;
  reg signed [16-1:0] __delay_data_2444__delay_2443__delay_2442___cond_2177;
  reg signed [16-1:0] __delay_data_2461__delay_2460__delay_2459___cond_2184;
  reg [16-1:0] __delay_data_2478__delay_2477__delay_2476___plus_2245;
  reg [1-1:0] __delay_data_2496__delay_2495__delay_2494__delay_2493___eq_2251;
  reg [1-1:0] __delay_data_2525__delay_2524__delay_2523__delay_2522___eq_2254;
  reg [1-1:0] __delay_data_2413__delay_2412__delay_2411____variable_2161;
  reg [16-1:0] __delay_data_2423__delay_2422__delay_2421___plus_2240;
  reg [13-1:0] __delay_data_2434__delay_2433__delay_2432____variable_2156;
  reg signed [16-1:0] __delay_data_2445__delay_2444__delay_2443___cond_2177;
  reg signed [16-1:0] __delay_data_2462__delay_2461__delay_2460___cond_2184;
  reg [16-1:0] __delay_data_2479__delay_2478__delay_2477___plus_2245;
  reg [1-1:0] __delay_data_2497__delay_2496__delay_2495__delay_2494___eq_2251;
  reg [1-1:0] __delay_data_2526__delay_2525__delay_2524__delay_2523___eq_2254;
  reg [1-1:0] __delay_data_2414__delay_2413__delay_2412____variable_2161;
  reg [16-1:0] __delay_data_2424__delay_2423__delay_2422___plus_2240;
  reg [13-1:0] __delay_data_2435__delay_2434__delay_2433____variable_2156;
  reg signed [16-1:0] __delay_data_2446__delay_2445__delay_2444___cond_2177;
  reg signed [16-1:0] __delay_data_2463__delay_2462__delay_2461___cond_2184;
  reg [16-1:0] __delay_data_2480__delay_2479__delay_2478___plus_2245;
  reg [1-1:0] __delay_data_2498__delay_2497__delay_2496__delay_2495___eq_2251;
  reg [1-1:0] __delay_data_2527__delay_2526__delay_2525__delay_2524___eq_2254;
  reg [1-1:0] __delay_data_2415__delay_2414__delay_2413____variable_2161;
  reg [16-1:0] __delay_data_2425__delay_2424__delay_2423___plus_2240;
  reg [13-1:0] __delay_data_2436__delay_2435__delay_2434____variable_2156;
  reg signed [16-1:0] __delay_data_2447__delay_2446__delay_2445___cond_2177;
  reg signed [16-1:0] __delay_data_2464__delay_2463__delay_2462___cond_2184;
  reg [16-1:0] __delay_data_2481__delay_2480__delay_2479___plus_2245;
  reg [1-1:0] __delay_data_2499__delay_2498__delay_2497__delay_2496___eq_2251;
  reg [1-1:0] __delay_data_2528__delay_2527__delay_2526__delay_2525___eq_2254;
  wire signed [32-1:0] __substreamoutput_data_2236;
  assign __substreamoutput_data_2236 = mul_18_z_data;
  reg signed [64-1:0] __variable_wdata_1302;
  assign add_tree_15_var0_data = __variable_wdata_1302;
  assign _add_tree_15_is_root = ((_stream_matmul_11_busy)? 0 : 1) && 1;
  assign _add_tree_15_stream_oready = ((_stream_matmul_11_busy)? _stream_matmul_11_stream_oready : 1) && _add_tree_15_stream_internal_oready;
  reg [1-1:0] __delay_data_2416__delay_2415__delay_2414____variable_2161;
  reg [16-1:0] __delay_data_2426__delay_2425__delay_2424___plus_2240;
  reg [13-1:0] __delay_data_2437__delay_2436__delay_2435____variable_2156;
  reg signed [16-1:0] __delay_data_2448__delay_2447__delay_2446___cond_2177;
  reg signed [16-1:0] __delay_data_2465__delay_2464__delay_2463___cond_2184;
  reg [16-1:0] __delay_data_2482__delay_2481__delay_2480___plus_2245;
  reg [1-1:0] __delay_data_2500__delay_2499__delay_2498__delay_2497___eq_2251;
  reg [1-1:0] __delay_data_2529__delay_2528__delay_2527__delay_2526___eq_2254;
  wire signed [64-1:0] __substreamoutput_data_2238;
  assign __substreamoutput_data_2238 = add_tree_15_sum_data;
  assign _acc_14_is_root = ((_stream_matmul_11_busy)? 0 : 1) && (((_stream_conv2d_4_busy)? 0 : 1) && 1);
  assign _acc_14_stream_oready = ((_stream_matmul_11_busy)? _stream_matmul_11_stream_oready : 1) && (((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _acc_14_stream_internal_oready);
  reg signed [16-1:0] __delay_data_2449__delay_2448__delay_2447___cond_2177;
  reg signed [16-1:0] __delay_data_2466__delay_2465__delay_2464___cond_2184;
  reg [16-1:0] __delay_data_2483__delay_2482__delay_2481___plus_2245;
  reg [1-1:0] __delay_data_2501__delay_2500__delay_2499__delay_2498___eq_2251;
  reg [1-1:0] __delay_data_2530__delay_2529__delay_2528__delay_2527___eq_2254;
  reg signed [16-1:0] __delay_data_2450__delay_2449__delay_2448___cond_2177;
  reg signed [16-1:0] __delay_data_2467__delay_2466__delay_2465___cond_2184;
  reg [16-1:0] __delay_data_2484__delay_2483__delay_2482___plus_2245;
  reg [1-1:0] __delay_data_2502__delay_2501__delay_2500__delay_2499___eq_2251;
  reg [1-1:0] __delay_data_2531__delay_2530__delay_2529__delay_2528___eq_2254;
  reg signed [16-1:0] __delay_data_2451__delay_2450__delay_2449___cond_2177;
  reg signed [16-1:0] __delay_data_2468__delay_2467__delay_2466___cond_2184;
  reg [16-1:0] __delay_data_2485__delay_2484__delay_2483___plus_2245;
  reg [1-1:0] __delay_data_2503__delay_2502__delay_2501__delay_2500___eq_2251;
  reg [1-1:0] __delay_data_2532__delay_2531__delay_2530__delay_2529___eq_2254;
  reg signed [16-1:0] __delay_data_2452__delay_2451__delay_2450___cond_2177;
  reg signed [16-1:0] __delay_data_2469__delay_2468__delay_2467___cond_2184;
  reg [16-1:0] __delay_data_2486__delay_2485__delay_2484___plus_2245;
  reg [1-1:0] __delay_data_2504__delay_2503__delay_2502__delay_2501___eq_2251;
  reg [1-1:0] __delay_data_2533__delay_2532__delay_2531__delay_2530___eq_2254;
  reg signed [16-1:0] __delay_data_2453__delay_2452__delay_2451___cond_2177;
  reg signed [16-1:0] __delay_data_2470__delay_2469__delay_2468___cond_2184;
  reg [16-1:0] __delay_data_2487__delay_2486__delay_2485___plus_2245;
  reg [1-1:0] __delay_data_2505__delay_2504__delay_2503__delay_2502___eq_2251;
  reg [1-1:0] __delay_data_2534__delay_2533__delay_2532__delay_2531___eq_2254;
  reg signed [16-1:0] __delay_data_2454__delay_2453__delay_2452___cond_2177;
  reg signed [16-1:0] __delay_data_2471__delay_2470__delay_2469___cond_2184;
  reg [16-1:0] __delay_data_2488__delay_2487__delay_2486___plus_2245;
  reg [1-1:0] __delay_data_2506__delay_2505__delay_2504__delay_2503___eq_2251;
  reg [1-1:0] __delay_data_2535__delay_2534__delay_2533__delay_2532___eq_2254;
  wire signed [64-1:0] __substreamoutput_data_2241;
  assign __substreamoutput_data_2241 = acc_14_sum_data;
  wire [1-1:0] __substreamoutput_data_2242;
  assign __substreamoutput_data_2242 = acc_14_valid_data;
  reg signed [64-1:0] _plus_data_2243;
  reg signed [16-1:0] __delay_data_2472__delay_2471__delay_2470___cond_2184;
  reg [16-1:0] __delay_data_2489__delay_2488__delay_2487___plus_2245;
  reg [1-1:0] __delay_data_2507__delay_2506__delay_2505__delay_2504___eq_2251;
  reg [1-1:0] __delay_data_2536__delay_2535__delay_2534__delay_2533___eq_2254;
  reg [1-1:0] __delay_data_2548__substreamoutput_2242;
  assign _mul_rshift_round_clip_17_is_root = ((_stream_matmul_11_busy)? 0 : 1) && (((_stream_conv2d_4_busy)? 0 : 1) && 1);
  assign _mul_rshift_round_clip_17_stream_oready = ((_stream_matmul_11_busy)? _stream_matmul_11_stream_oready : 1) && (((_stream_conv2d_4_busy)? _stream_conv2d_4_stream_oready : 1) && _mul_rshift_round_clip_17_stream_internal_oready);
  assign _stream_matmul_11_stream_internal_oready = ((_stream_matmul_11_busy)? _mul_rshift_round_clip_17_stream_internal_oready : 1) && (((_stream_matmul_11_busy)? _acc_14_stream_internal_oready : 1) && (((_stream_matmul_11_busy)? _add_tree_15_stream_internal_oready : 1) && (((_stream_matmul_11_busy)? _mul_18_stream_internal_oready : 1) && 1)));
  reg [1-1:0] __delay_data_2508__delay_2507__delay_2506__delay_2505___eq_2251;
  reg [1-1:0] __delay_data_2537__delay_2536__delay_2535__delay_2534___eq_2254;
  reg [1-1:0] __delay_data_2549__delay_2548__substreamoutput_2242;
  reg [1-1:0] __delay_data_2509__delay_2508__delay_2507__delay_2506___eq_2251;
  reg [1-1:0] __delay_data_2538__delay_2537__delay_2536__delay_2535___eq_2254;
  reg [1-1:0] __delay_data_2550__delay_2549____substreamoutput_2242;
  reg [1-1:0] __delay_data_2510__delay_2509__delay_2508__delay_2507___eq_2251;
  reg [1-1:0] __delay_data_2539__delay_2538__delay_2537__delay_2536___eq_2254;
  reg [1-1:0] __delay_data_2551__delay_2550____substreamoutput_2242;
  reg [1-1:0] __delay_data_2511__delay_2510__delay_2509__delay_2508___eq_2251;
  reg [1-1:0] __delay_data_2540__delay_2539__delay_2538__delay_2537___eq_2254;
  reg [1-1:0] __delay_data_2552__delay_2551____substreamoutput_2242;
  reg [1-1:0] __delay_data_2512__delay_2511__delay_2510__delay_2509___eq_2251;
  reg [1-1:0] __delay_data_2541__delay_2540__delay_2539__delay_2538___eq_2254;
  reg [1-1:0] __delay_data_2553__delay_2552____substreamoutput_2242;
  reg [1-1:0] __delay_data_2513__delay_2512__delay_2511__delay_2510___eq_2251;
  reg [1-1:0] __delay_data_2542__delay_2541__delay_2540__delay_2539___eq_2254;
  reg [1-1:0] __delay_data_2554__delay_2553____substreamoutput_2242;
  reg [1-1:0] __delay_data_2514__delay_2513__delay_2512__delay_2511___eq_2251;
  reg [1-1:0] __delay_data_2543__delay_2542__delay_2541__delay_2540___eq_2254;
  reg [1-1:0] __delay_data_2555__delay_2554____substreamoutput_2242;
  reg [1-1:0] __delay_data_2515__delay_2514__delay_2513__delay_2512___eq_2251;
  reg [1-1:0] __delay_data_2544__delay_2543__delay_2542__delay_2541___eq_2254;
  reg [1-1:0] __delay_data_2556__delay_2555____substreamoutput_2242;
  reg [1-1:0] __delay_data_2516__delay_2515__delay_2514__delay_2513___eq_2251;
  reg [1-1:0] __delay_data_2545__delay_2544__delay_2543__delay_2542___eq_2254;
  reg [1-1:0] __delay_data_2557__delay_2556____substreamoutput_2242;
  wire signed [16-1:0] __substreamoutput_data_2246;
  assign __substreamoutput_data_2246 = mul_rshift_round_clip_17_z_data;
  reg [1-1:0] _greaterthan_data_2248;
  reg signed [16-1:0] __delay_data_2490__substreamoutput_2246;
  reg [1-1:0] __delay_data_2517__delay_2516__delay_2515__delay_2514___eq_2251;
  reg [1-1:0] __delay_data_2546__delay_2545__delay_2544__delay_2543___eq_2254;
  reg [1-1:0] __delay_data_2558__delay_2557____substreamoutput_2242;
  reg signed [16-1:0] _cond_data_2250;
  reg [1-1:0] __delay_data_2518__delay_2517__delay_2516__delay_2515___eq_2251;
  reg signed [16-1:0] __delay_data_2519__delay_2490__substreamoutput_2246;
  reg [1-1:0] __delay_data_2547__delay_2546__delay_2545__delay_2544___eq_2254;
  reg [1-1:0] __delay_data_2559__delay_2558____substreamoutput_2242;
  wire signed [16-1:0] _cond_data_2253;
  assign _cond_data_2253 = (__delay_data_2518__delay_2517__delay_2516__delay_2515___eq_2251)? _cond_data_2250 : __delay_data_2519__delay_2490__substreamoutput_2246;
  wire signed [16-1:0] _cond_data_2256;
  assign _cond_data_2256 = (__delay_data_2547__delay_2546__delay_2545__delay_2544___eq_2254)? __delay_data_2519__delay_2490__substreamoutput_2246 : _cond_data_2253;
  wire signed [16-1:0] _reinterpretcast_src_2257;
  assign _reinterpretcast_src_2257 = _cond_data_2256;
  wire signed [16-1:0] _reinterpretcast_data_2257;
  assign _reinterpretcast_data_2257 = _reinterpretcast_src_2257;
  wire signed [16-1:0] stream_matmul_11_sink_26_data;
  assign stream_matmul_11_sink_26_data = _reinterpretcast_data_2257;
  wire [1-1:0] stream_matmul_11_sink_27_data;
  assign stream_matmul_11_sink_27_data = __delay_data_2559__delay_2558____substreamoutput_2242;
  wire _set_flag_1356;
  assign _set_flag_1356 = matmul_11_comp_fsm == 3;
  reg [13-1:0] __variable_wdata_2156;
  assign stream_matmul_11_parameter_0_data = __variable_wdata_2156;
  wire _set_flag_1357;
  assign _set_flag_1357 = matmul_11_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_2157;
  assign stream_matmul_11_parameter_1_data = __variable_wdata_2157;
  wire _set_flag_1358;
  assign _set_flag_1358 = matmul_11_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_2158;
  assign stream_matmul_11_parameter_2_data = __variable_wdata_2158;
  wire _set_flag_1359;
  assign _set_flag_1359 = matmul_11_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_2159;
  assign stream_matmul_11_parameter_3_data = __variable_wdata_2159;
  wire _set_flag_1360;
  assign _set_flag_1360 = matmul_11_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_2160;
  assign stream_matmul_11_parameter_4_data = __variable_wdata_2160;
  wire _set_flag_1361;
  assign _set_flag_1361 = matmul_11_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_2171;
  assign stream_matmul_11_parameter_6_data = __variable_wdata_2171;
  reg [32-1:0] _source_stream_matmul_11_source_7_pat_cur_offset_0;
  reg [32-1:0] _source_stream_matmul_11_source_7_pat_cur_offset_1;
  reg [32-1:0] _source_stream_matmul_11_source_7_pat_cur_offset_2;
  reg [32-1:0] _source_stream_matmul_11_source_7_pat_cur_offset_3;
  reg [33-1:0] _source_stream_matmul_11_source_7_pat_size_0;
  reg [33-1:0] _source_stream_matmul_11_source_7_pat_size_1;
  reg [33-1:0] _source_stream_matmul_11_source_7_pat_size_2;
  reg [33-1:0] _source_stream_matmul_11_source_7_pat_size_3;
  reg [32-1:0] _source_stream_matmul_11_source_7_pat_stride_0;
  reg [32-1:0] _source_stream_matmul_11_source_7_pat_stride_1;
  reg [32-1:0] _source_stream_matmul_11_source_7_pat_stride_2;
  reg [32-1:0] _source_stream_matmul_11_source_7_pat_stride_3;
  reg [33-1:0] _source_stream_matmul_11_source_7_pat_count_0;
  reg [33-1:0] _source_stream_matmul_11_source_7_pat_count_1;
  reg [33-1:0] _source_stream_matmul_11_source_7_pat_count_2;
  reg [33-1:0] _source_stream_matmul_11_source_7_pat_count_3;
  reg [33-1:0] _source_stream_matmul_11_source_7_pat_size_buf_0;
  reg [33-1:0] _source_stream_matmul_11_source_7_pat_size_buf_1;
  reg [33-1:0] _source_stream_matmul_11_source_7_pat_size_buf_2;
  reg [33-1:0] _source_stream_matmul_11_source_7_pat_size_buf_3;
  reg [32-1:0] _source_stream_matmul_11_source_7_pat_stride_buf_0;
  reg [32-1:0] _source_stream_matmul_11_source_7_pat_stride_buf_1;
  reg [32-1:0] _source_stream_matmul_11_source_7_pat_stride_buf_2;
  reg [32-1:0] _source_stream_matmul_11_source_7_pat_stride_buf_3;
  wire _set_flag_1362;
  assign _set_flag_1362 = matmul_11_comp_fsm == 3;
  wire [1-1:0] read_rtl_bank_1363;
  assign read_rtl_bank_1363 = _stream_matmul_11_source_7_source_ram_raddr;
  reg [1-1:0] _tmp_1364;
  assign ram_w16_l512_id1_0_0_addr = (_stream_matmul_11_stream_oready && _stream_matmul_11_source_7_source_ram_renable && (_stream_matmul_11_source_7_source_sel == 1))? _stream_matmul_11_source_7_source_ram_raddr >> 1 : 
                                     (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_30_source_ram_renable && (_stream_conv2d_4_source_30_source_sel == 13))? _stream_conv2d_4_source_30_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id1_0_0_enable = (_stream_matmul_11_stream_oready && _stream_matmul_11_source_7_source_ram_renable && (_stream_matmul_11_source_7_source_sel == 1))? 1'd1 : 
                                       (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_30_source_ram_renable && (_stream_conv2d_4_source_30_source_sel == 13))? 1'd1 : 0;
  localparam _tmp_1365 = 1;
  wire [_tmp_1365-1:0] _tmp_1366;
  assign _tmp_1366 = _stream_matmul_11_stream_oready && _stream_matmul_11_source_7_source_ram_renable && (_stream_matmul_11_source_7_source_sel == 1);
  reg [_tmp_1365-1:0] __tmp_1366_1;
  assign ram_w16_l512_id1_1_0_addr = (_stream_matmul_11_stream_oready && _stream_matmul_11_source_7_source_ram_renable && (_stream_matmul_11_source_7_source_sel == 1))? _stream_matmul_11_source_7_source_ram_raddr >> 1 : 
                                     (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_30_source_ram_renable && (_stream_conv2d_4_source_30_source_sel == 13))? _stream_conv2d_4_source_30_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id1_1_0_enable = (_stream_matmul_11_stream_oready && _stream_matmul_11_source_7_source_ram_renable && (_stream_matmul_11_source_7_source_sel == 1))? 1'd1 : 
                                       (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_30_source_ram_renable && (_stream_conv2d_4_source_30_source_sel == 13))? 1'd1 : 0;
  localparam _tmp_1367 = 1;
  wire [_tmp_1367-1:0] _tmp_1368;
  assign _tmp_1368 = _stream_matmul_11_stream_oready && _stream_matmul_11_source_7_source_ram_renable && (_stream_matmul_11_source_7_source_sel == 1);
  reg [_tmp_1367-1:0] __tmp_1368_1;
  wire signed [16-1:0] read_rtl_rdata_1369;
  wire read_rtl_rvalid_1370;
  assign read_rtl_rdata_1369 = (_tmp_1364 == 0)? ram_w16_l512_id1_0_0_rdata : 
                               (_tmp_1364 == 1)? ram_w16_l512_id1_1_0_rdata : 0;
  assign read_rtl_rvalid_1370 = __tmp_1366_1;
  assign _stream_matmul_11_source_7_source_ram_rdata = (_stream_matmul_11_source_7_source_sel == 1)? read_rtl_rdata_1369 : 'hx;
  reg [16-1:0] __variable_wdata_2172;
  assign stream_matmul_11_source_7_data = __variable_wdata_2172;
  reg [32-1:0] _stream_matmul_11_source_7_source_pat_fsm_0;
  localparam _stream_matmul_11_source_7_source_pat_fsm_0_init = 0;
  wire [32-1:0] _stream_matmul_11_source_7_source_pat_all_offset;
  assign _stream_matmul_11_source_7_source_pat_all_offset = _stream_matmul_11_source_7_source_offset_buf + _source_stream_matmul_11_source_7_pat_cur_offset_0 + _source_stream_matmul_11_source_7_pat_cur_offset_1 + _source_stream_matmul_11_source_7_pat_cur_offset_2 + _source_stream_matmul_11_source_7_pat_cur_offset_3;
  wire _set_flag_1371;
  assign _set_flag_1371 = matmul_11_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_2178;
  assign stream_matmul_11_parameter_8_data = __variable_wdata_2178;
  reg [32-1:0] _source_stream_matmul_11_source_9_pat_cur_offset_0;
  reg [32-1:0] _source_stream_matmul_11_source_9_pat_cur_offset_1;
  reg [32-1:0] _source_stream_matmul_11_source_9_pat_cur_offset_2;
  reg [32-1:0] _source_stream_matmul_11_source_9_pat_cur_offset_3;
  reg [33-1:0] _source_stream_matmul_11_source_9_pat_size_0;
  reg [33-1:0] _source_stream_matmul_11_source_9_pat_size_1;
  reg [33-1:0] _source_stream_matmul_11_source_9_pat_size_2;
  reg [33-1:0] _source_stream_matmul_11_source_9_pat_size_3;
  reg [32-1:0] _source_stream_matmul_11_source_9_pat_stride_0;
  reg [32-1:0] _source_stream_matmul_11_source_9_pat_stride_1;
  reg [32-1:0] _source_stream_matmul_11_source_9_pat_stride_2;
  reg [32-1:0] _source_stream_matmul_11_source_9_pat_stride_3;
  reg [33-1:0] _source_stream_matmul_11_source_9_pat_count_0;
  reg [33-1:0] _source_stream_matmul_11_source_9_pat_count_1;
  reg [33-1:0] _source_stream_matmul_11_source_9_pat_count_2;
  reg [33-1:0] _source_stream_matmul_11_source_9_pat_count_3;
  reg [33-1:0] _source_stream_matmul_11_source_9_pat_size_buf_0;
  reg [33-1:0] _source_stream_matmul_11_source_9_pat_size_buf_1;
  reg [33-1:0] _source_stream_matmul_11_source_9_pat_size_buf_2;
  reg [33-1:0] _source_stream_matmul_11_source_9_pat_size_buf_3;
  reg [32-1:0] _source_stream_matmul_11_source_9_pat_stride_buf_0;
  reg [32-1:0] _source_stream_matmul_11_source_9_pat_stride_buf_1;
  reg [32-1:0] _source_stream_matmul_11_source_9_pat_stride_buf_2;
  reg [32-1:0] _source_stream_matmul_11_source_9_pat_stride_buf_3;
  wire _set_flag_1372;
  assign _set_flag_1372 = matmul_11_comp_fsm == 3;
  wire [1-1:0] read_rtl_bank_1373;
  assign read_rtl_bank_1373 = _stream_matmul_11_source_9_source_ram_raddr;
  reg [1-1:0] _tmp_1374;
  assign ram_w16_l512_id2_0_0_addr = (_stream_matmul_11_stream_oready && _stream_matmul_11_source_9_source_ram_renable && (_stream_matmul_11_source_9_source_sel == 2))? _stream_matmul_11_source_9_source_ram_raddr >> 1 : 
                                     (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_31_source_ram_renable && (_stream_conv2d_4_source_31_source_sel == 14))? _stream_conv2d_4_source_31_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id2_0_0_enable = (_stream_matmul_11_stream_oready && _stream_matmul_11_source_9_source_ram_renable && (_stream_matmul_11_source_9_source_sel == 2))? 1'd1 : 
                                       (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_31_source_ram_renable && (_stream_conv2d_4_source_31_source_sel == 14))? 1'd1 : 0;
  localparam _tmp_1375 = 1;
  wire [_tmp_1375-1:0] _tmp_1376;
  assign _tmp_1376 = _stream_matmul_11_stream_oready && _stream_matmul_11_source_9_source_ram_renable && (_stream_matmul_11_source_9_source_sel == 2);
  reg [_tmp_1375-1:0] __tmp_1376_1;
  assign ram_w16_l512_id2_1_0_addr = (_stream_matmul_11_stream_oready && _stream_matmul_11_source_9_source_ram_renable && (_stream_matmul_11_source_9_source_sel == 2))? _stream_matmul_11_source_9_source_ram_raddr >> 1 : 
                                     (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_31_source_ram_renable && (_stream_conv2d_4_source_31_source_sel == 14))? _stream_conv2d_4_source_31_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id2_1_0_enable = (_stream_matmul_11_stream_oready && _stream_matmul_11_source_9_source_ram_renable && (_stream_matmul_11_source_9_source_sel == 2))? 1'd1 : 
                                       (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_31_source_ram_renable && (_stream_conv2d_4_source_31_source_sel == 14))? 1'd1 : 0;
  localparam _tmp_1377 = 1;
  wire [_tmp_1377-1:0] _tmp_1378;
  assign _tmp_1378 = _stream_matmul_11_stream_oready && _stream_matmul_11_source_9_source_ram_renable && (_stream_matmul_11_source_9_source_sel == 2);
  reg [_tmp_1377-1:0] __tmp_1378_1;
  wire signed [16-1:0] read_rtl_rdata_1379;
  wire read_rtl_rvalid_1380;
  assign read_rtl_rdata_1379 = (_tmp_1374 == 0)? ram_w16_l512_id2_0_0_rdata : 
                               (_tmp_1374 == 1)? ram_w16_l512_id2_1_0_rdata : 0;
  assign read_rtl_rvalid_1380 = __tmp_1376_1;
  assign _stream_matmul_11_source_9_source_ram_rdata = (_stream_matmul_11_source_9_source_sel == 2)? read_rtl_rdata_1379 : 'hx;
  reg [16-1:0] __variable_wdata_2179;
  assign stream_matmul_11_source_9_data = __variable_wdata_2179;
  reg [32-1:0] _stream_matmul_11_source_9_source_pat_fsm_1;
  localparam _stream_matmul_11_source_9_source_pat_fsm_1_init = 0;
  wire [32-1:0] _stream_matmul_11_source_9_source_pat_all_offset;
  assign _stream_matmul_11_source_9_source_pat_all_offset = _stream_matmul_11_source_9_source_offset_buf + _source_stream_matmul_11_source_9_pat_cur_offset_0 + _source_stream_matmul_11_source_9_pat_cur_offset_1 + _source_stream_matmul_11_source_9_pat_cur_offset_2 + _source_stream_matmul_11_source_9_pat_cur_offset_3;
  wire _set_flag_1381;
  assign _set_flag_1381 = matmul_11_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_2185;
  assign stream_matmul_11_parameter_10_data = __variable_wdata_2185;
  wire _set_flag_1382;
  assign _set_flag_1382 = matmul_11_comp_fsm == 3;
  reg [16-1:0] __variable_wdata_2186;
  assign stream_matmul_11_source_11_data = __variable_wdata_2186;
  wire _set_flag_1383;
  assign _set_flag_1383 = matmul_11_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_2192;
  assign stream_matmul_11_parameter_12_data = __variable_wdata_2192;
  wire _set_flag_1384;
  assign _set_flag_1384 = matmul_11_comp_fsm == 3;
  reg [16-1:0] __variable_wdata_2193;
  assign stream_matmul_11_source_13_data = __variable_wdata_2193;
  wire _set_flag_1385;
  assign _set_flag_1385 = matmul_11_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_2199;
  assign stream_matmul_11_parameter_14_data = __variable_wdata_2199;
  wire _set_flag_1386;
  assign _set_flag_1386 = matmul_11_comp_fsm == 3;
  reg [16-1:0] __variable_wdata_2200;
  assign stream_matmul_11_source_15_data = __variable_wdata_2200;
  wire _set_flag_1387;
  assign _set_flag_1387 = matmul_11_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_2206;
  assign stream_matmul_11_parameter_16_data = __variable_wdata_2206;
  wire _set_flag_1388;
  assign _set_flag_1388 = matmul_11_comp_fsm == 3;
  reg [1-1:0] __variable_wdata_2207;
  assign stream_matmul_11_parameter_17_data = __variable_wdata_2207;
  wire _set_flag_1389;
  assign _set_flag_1389 = matmul_11_comp_fsm == 3;
  reg [5-1:0] __variable_wdata_2208;
  assign stream_matmul_11_parameter_18_data = __variable_wdata_2208;
  wire _set_flag_1390;
  assign _set_flag_1390 = matmul_11_comp_fsm == 3;
  reg [2-1:0] __variable_wdata_2209;
  assign stream_matmul_11_parameter_19_data = __variable_wdata_2209;
  reg [32-1:0] _source_stream_matmul_11_source_20_pat_cur_offset_0;
  reg [32-1:0] _source_stream_matmul_11_source_20_pat_cur_offset_1;
  reg [32-1:0] _source_stream_matmul_11_source_20_pat_cur_offset_2;
  reg [32-1:0] _source_stream_matmul_11_source_20_pat_cur_offset_3;
  reg [33-1:0] _source_stream_matmul_11_source_20_pat_size_0;
  reg [33-1:0] _source_stream_matmul_11_source_20_pat_size_1;
  reg [33-1:0] _source_stream_matmul_11_source_20_pat_size_2;
  reg [33-1:0] _source_stream_matmul_11_source_20_pat_size_3;
  reg [32-1:0] _source_stream_matmul_11_source_20_pat_stride_0;
  reg [32-1:0] _source_stream_matmul_11_source_20_pat_stride_1;
  reg [32-1:0] _source_stream_matmul_11_source_20_pat_stride_2;
  reg [32-1:0] _source_stream_matmul_11_source_20_pat_stride_3;
  reg [33-1:0] _source_stream_matmul_11_source_20_pat_count_0;
  reg [33-1:0] _source_stream_matmul_11_source_20_pat_count_1;
  reg [33-1:0] _source_stream_matmul_11_source_20_pat_count_2;
  reg [33-1:0] _source_stream_matmul_11_source_20_pat_count_3;
  reg [33-1:0] _source_stream_matmul_11_source_20_pat_size_buf_0;
  reg [33-1:0] _source_stream_matmul_11_source_20_pat_size_buf_1;
  reg [33-1:0] _source_stream_matmul_11_source_20_pat_size_buf_2;
  reg [33-1:0] _source_stream_matmul_11_source_20_pat_size_buf_3;
  reg [32-1:0] _source_stream_matmul_11_source_20_pat_stride_buf_0;
  reg [32-1:0] _source_stream_matmul_11_source_20_pat_stride_buf_1;
  reg [32-1:0] _source_stream_matmul_11_source_20_pat_stride_buf_2;
  reg [32-1:0] _source_stream_matmul_11_source_20_pat_stride_buf_3;
  wire _set_flag_1391;
  assign _set_flag_1391 = matmul_11_comp_fsm == 3;
  wire [1-1:0] read_rtl_bank_1392;
  assign read_rtl_bank_1392 = _stream_matmul_11_source_20_source_ram_raddr;
  reg [1-1:0] _tmp_1393;
  assign ram_w16_l8192_id0_0_0_addr = (_stream_matmul_11_stream_oready && _stream_matmul_11_source_20_source_ram_renable && (_stream_matmul_11_source_20_source_sel == 3))? _stream_matmul_11_source_20_source_ram_raddr >> 1 : 
                                      (_stream_max_pool_serial_6_stream_oready && _stream_max_pool_serial_6_sink_5_sink_wenable && (_stream_max_pool_serial_6_sink_5_sink_sel == 2) && (write_rtl_bank_1233 == 0))? _stream_max_pool_serial_6_sink_5_sink_waddr >> 1 : 'hx;
  assign ram_w16_l8192_id0_0_0_enable = (_stream_matmul_11_stream_oready && _stream_matmul_11_source_20_source_ram_renable && (_stream_matmul_11_source_20_source_sel == 3))? 1'd1 : 
                                        (_stream_max_pool_serial_6_stream_oready && _stream_max_pool_serial_6_sink_5_sink_wenable && (_stream_max_pool_serial_6_sink_5_sink_sel == 2) && (write_rtl_bank_1233 == 0))? 1'd1 : 0;
  localparam _tmp_1394 = 1;
  wire [_tmp_1394-1:0] _tmp_1395;
  assign _tmp_1395 = _stream_matmul_11_stream_oready && _stream_matmul_11_source_20_source_ram_renable && (_stream_matmul_11_source_20_source_sel == 3);
  reg [_tmp_1394-1:0] __tmp_1395_1;
  assign ram_w16_l8192_id0_1_0_addr = (_stream_matmul_11_stream_oready && _stream_matmul_11_source_20_source_ram_renable && (_stream_matmul_11_source_20_source_sel == 3))? _stream_matmul_11_source_20_source_ram_raddr >> 1 : 
                                      (_stream_max_pool_serial_6_stream_oready && _stream_max_pool_serial_6_sink_5_sink_wenable && (_stream_max_pool_serial_6_sink_5_sink_sel == 2) && (write_rtl_bank_1233 == 1))? _stream_max_pool_serial_6_sink_5_sink_waddr >> 1 : 'hx;
  assign ram_w16_l8192_id0_1_0_enable = (_stream_matmul_11_stream_oready && _stream_matmul_11_source_20_source_ram_renable && (_stream_matmul_11_source_20_source_sel == 3))? 1'd1 : 
                                        (_stream_max_pool_serial_6_stream_oready && _stream_max_pool_serial_6_sink_5_sink_wenable && (_stream_max_pool_serial_6_sink_5_sink_sel == 2) && (write_rtl_bank_1233 == 1))? 1'd1 : 0;
  localparam _tmp_1396 = 1;
  wire [_tmp_1396-1:0] _tmp_1397;
  assign _tmp_1397 = _stream_matmul_11_stream_oready && _stream_matmul_11_source_20_source_ram_renable && (_stream_matmul_11_source_20_source_sel == 3);
  reg [_tmp_1396-1:0] __tmp_1397_1;
  wire signed [16-1:0] read_rtl_rdata_1398;
  wire read_rtl_rvalid_1399;
  assign read_rtl_rdata_1398 = (_tmp_1393 == 0)? ram_w16_l8192_id0_0_0_rdata : 
                               (_tmp_1393 == 1)? ram_w16_l8192_id0_1_0_rdata : 0;
  assign read_rtl_rvalid_1399 = __tmp_1395_1;
  assign _stream_matmul_11_source_20_source_ram_rdata = (_stream_matmul_11_source_20_source_sel == 3)? read_rtl_rdata_1398 : 'hx;
  reg [16-1:0] __variable_wdata_2210;
  assign stream_matmul_11_source_20_data = __variable_wdata_2210;
  reg [32-1:0] _stream_matmul_11_source_20_source_pat_fsm_2;
  localparam _stream_matmul_11_source_20_source_pat_fsm_2_init = 0;
  wire [32-1:0] _stream_matmul_11_source_20_source_pat_all_offset;
  assign _stream_matmul_11_source_20_source_pat_all_offset = _stream_matmul_11_source_20_source_offset_buf + _source_stream_matmul_11_source_20_pat_cur_offset_0 + _source_stream_matmul_11_source_20_pat_cur_offset_1 + _source_stream_matmul_11_source_20_pat_cur_offset_2 + _source_stream_matmul_11_source_20_pat_cur_offset_3;
  reg [32-1:0] _source_stream_matmul_11_source_21_pat_cur_offset_0;
  reg [32-1:0] _source_stream_matmul_11_source_21_pat_cur_offset_1;
  reg [32-1:0] _source_stream_matmul_11_source_21_pat_cur_offset_2;
  reg [32-1:0] _source_stream_matmul_11_source_21_pat_cur_offset_3;
  reg [33-1:0] _source_stream_matmul_11_source_21_pat_size_0;
  reg [33-1:0] _source_stream_matmul_11_source_21_pat_size_1;
  reg [33-1:0] _source_stream_matmul_11_source_21_pat_size_2;
  reg [33-1:0] _source_stream_matmul_11_source_21_pat_size_3;
  reg [32-1:0] _source_stream_matmul_11_source_21_pat_stride_0;
  reg [32-1:0] _source_stream_matmul_11_source_21_pat_stride_1;
  reg [32-1:0] _source_stream_matmul_11_source_21_pat_stride_2;
  reg [32-1:0] _source_stream_matmul_11_source_21_pat_stride_3;
  reg [33-1:0] _source_stream_matmul_11_source_21_pat_count_0;
  reg [33-1:0] _source_stream_matmul_11_source_21_pat_count_1;
  reg [33-1:0] _source_stream_matmul_11_source_21_pat_count_2;
  reg [33-1:0] _source_stream_matmul_11_source_21_pat_count_3;
  reg [33-1:0] _source_stream_matmul_11_source_21_pat_size_buf_0;
  reg [33-1:0] _source_stream_matmul_11_source_21_pat_size_buf_1;
  reg [33-1:0] _source_stream_matmul_11_source_21_pat_size_buf_2;
  reg [33-1:0] _source_stream_matmul_11_source_21_pat_size_buf_3;
  reg [32-1:0] _source_stream_matmul_11_source_21_pat_stride_buf_0;
  reg [32-1:0] _source_stream_matmul_11_source_21_pat_stride_buf_1;
  reg [32-1:0] _source_stream_matmul_11_source_21_pat_stride_buf_2;
  reg [32-1:0] _source_stream_matmul_11_source_21_pat_stride_buf_3;
  wire _set_flag_1400;
  assign _set_flag_1400 = matmul_11_comp_fsm == 3;
  wire [1-1:0] read_rtl_bank_1401;
  assign read_rtl_bank_1401 = _stream_matmul_11_source_21_source_ram_raddr;
  reg [1-1:0] _tmp_1402;
  assign ram_w16_l32768_id0_0_0_addr = (_stream_matmul_11_stream_oready && _stream_matmul_11_source_21_source_ram_renable && (_stream_matmul_11_source_21_source_sel == 4))? _stream_matmul_11_source_21_source_ram_raddr >> 1 : 
                                       (_stream_max_pool_serial_6_stream_oready && _stream_max_pool_serial_6_source_1_source_ram_renable && (_stream_max_pool_serial_6_source_1_source_sel == 1))? _stream_max_pool_serial_6_source_1_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l32768_id0_0_0_enable = (_stream_matmul_11_stream_oready && _stream_matmul_11_source_21_source_ram_renable && (_stream_matmul_11_source_21_source_sel == 4))? 1'd1 : 
                                         (_stream_max_pool_serial_6_stream_oready && _stream_max_pool_serial_6_source_1_source_ram_renable && (_stream_max_pool_serial_6_source_1_source_sel == 1))? 1'd1 : 0;
  localparam _tmp_1403 = 1;
  wire [_tmp_1403-1:0] _tmp_1404;
  assign _tmp_1404 = _stream_matmul_11_stream_oready && _stream_matmul_11_source_21_source_ram_renable && (_stream_matmul_11_source_21_source_sel == 4);
  reg [_tmp_1403-1:0] __tmp_1404_1;
  assign ram_w16_l32768_id0_1_0_addr = (_stream_matmul_11_stream_oready && _stream_matmul_11_source_21_source_ram_renable && (_stream_matmul_11_source_21_source_sel == 4))? _stream_matmul_11_source_21_source_ram_raddr >> 1 : 
                                       (_stream_max_pool_serial_6_stream_oready && _stream_max_pool_serial_6_source_1_source_ram_renable && (_stream_max_pool_serial_6_source_1_source_sel == 1))? _stream_max_pool_serial_6_source_1_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l32768_id0_1_0_enable = (_stream_matmul_11_stream_oready && _stream_matmul_11_source_21_source_ram_renable && (_stream_matmul_11_source_21_source_sel == 4))? 1'd1 : 
                                         (_stream_max_pool_serial_6_stream_oready && _stream_max_pool_serial_6_source_1_source_ram_renable && (_stream_max_pool_serial_6_source_1_source_sel == 1))? 1'd1 : 0;
  localparam _tmp_1405 = 1;
  wire [_tmp_1405-1:0] _tmp_1406;
  assign _tmp_1406 = _stream_matmul_11_stream_oready && _stream_matmul_11_source_21_source_ram_renable && (_stream_matmul_11_source_21_source_sel == 4);
  reg [_tmp_1405-1:0] __tmp_1406_1;
  wire signed [16-1:0] read_rtl_rdata_1407;
  wire read_rtl_rvalid_1408;
  assign read_rtl_rdata_1407 = (_tmp_1402 == 0)? ram_w16_l32768_id0_0_0_rdata : 
                               (_tmp_1402 == 1)? ram_w16_l32768_id0_1_0_rdata : 0;
  assign read_rtl_rvalid_1408 = __tmp_1404_1;
  assign _stream_matmul_11_source_21_source_ram_rdata = (_stream_matmul_11_source_21_source_sel == 4)? read_rtl_rdata_1407 : 'hx;
  reg [16-1:0] __variable_wdata_2224;
  assign stream_matmul_11_source_21_data = __variable_wdata_2224;
  reg [32-1:0] _stream_matmul_11_source_21_source_pat_fsm_3;
  localparam _stream_matmul_11_source_21_source_pat_fsm_3_init = 0;
  wire [32-1:0] _stream_matmul_11_source_21_source_pat_all_offset;
  assign _stream_matmul_11_source_21_source_pat_all_offset = _stream_matmul_11_source_21_source_offset_buf + _source_stream_matmul_11_source_21_pat_cur_offset_0 + _source_stream_matmul_11_source_21_pat_cur_offset_1 + _source_stream_matmul_11_source_21_pat_cur_offset_2 + _source_stream_matmul_11_source_21_pat_cur_offset_3;
  wire _set_flag_1409;
  assign _set_flag_1409 = matmul_11_comp_fsm == 3;
  reg _tmp_1410;
  reg _tmp_1411;
  reg _tmp_1412;
  reg _tmp_1413;
  reg _tmp_1414;
  reg _tmp_1415;
  reg _tmp_1416;
  reg _tmp_1417;
  reg _tmp_1418;
  reg _tmp_1419;
  reg _tmp_1420;
  reg _tmp_1421;
  reg _tmp_1422;
  reg _tmp_1423;
  reg _tmp_1424;
  reg _tmp_1425;
  reg _tmp_1426;
  reg _tmp_1427;
  reg _tmp_1428;
  reg _tmp_1429;
  reg _tmp_1430;
  reg _tmp_1431;
  reg _tmp_1432;
  reg _tmp_1433;
  reg _tmp_1434;
  reg _tmp_1435;
  reg _tmp_1436;
  reg _tmp_1437;
  reg _tmp_1438;
  reg _tmp_1439;
  reg _tmp_1440;
  localparam _tmp_1441 = 33;
  wire [_tmp_1441-1:0] _tmp_1442;
  assign _tmp_1442 = matmul_11_stream_out_local + matmul_11_out_page_comp_offset_buf;
  reg [_tmp_1441-1:0] _tmp_1443;
  reg [_tmp_1441-1:0] _tmp_1444;
  reg [_tmp_1441-1:0] _tmp_1445;
  reg [_tmp_1441-1:0] _tmp_1446;
  reg [_tmp_1441-1:0] _tmp_1447;
  reg [_tmp_1441-1:0] _tmp_1448;
  reg [_tmp_1441-1:0] _tmp_1449;
  reg [_tmp_1441-1:0] _tmp_1450;
  reg [_tmp_1441-1:0] _tmp_1451;
  reg [_tmp_1441-1:0] _tmp_1452;
  reg [_tmp_1441-1:0] _tmp_1453;
  reg [_tmp_1441-1:0] _tmp_1454;
  reg [_tmp_1441-1:0] _tmp_1455;
  reg [_tmp_1441-1:0] _tmp_1456;
  reg [_tmp_1441-1:0] _tmp_1457;
  reg [_tmp_1441-1:0] _tmp_1458;
  reg [_tmp_1441-1:0] _tmp_1459;
  reg [_tmp_1441-1:0] _tmp_1460;
  reg [_tmp_1441-1:0] _tmp_1461;
  reg [_tmp_1441-1:0] _tmp_1462;
  reg [_tmp_1441-1:0] _tmp_1463;
  reg [_tmp_1441-1:0] _tmp_1464;
  reg [_tmp_1441-1:0] _tmp_1465;
  reg [_tmp_1441-1:0] _tmp_1466;
  reg [_tmp_1441-1:0] _tmp_1467;
  reg [_tmp_1441-1:0] _tmp_1468;
  reg [_tmp_1441-1:0] _tmp_1469;
  reg [_tmp_1441-1:0] _tmp_1470;
  reg [_tmp_1441-1:0] _tmp_1471;
  reg [_tmp_1441-1:0] _tmp_1472;
  reg [_tmp_1441-1:0] _tmp_1473;
  reg [32-1:0] _tmp_1474;
  reg [32-1:0] _tmp_1475;
  reg [32-1:0] _tmp_1476;
  reg [32-1:0] _tmp_1477;
  reg [32-1:0] _tmp_1478;
  reg [32-1:0] _tmp_1479;
  reg [32-1:0] _tmp_1480;
  reg [32-1:0] _tmp_1481;
  reg [32-1:0] _tmp_1482;
  reg [32-1:0] _tmp_1483;
  reg [32-1:0] _tmp_1484;
  reg [32-1:0] _tmp_1485;
  reg [32-1:0] _tmp_1486;
  reg [32-1:0] _tmp_1487;
  reg [32-1:0] _tmp_1488;
  reg [32-1:0] _tmp_1489;
  reg [32-1:0] _tmp_1490;
  reg [32-1:0] _tmp_1491;
  reg [32-1:0] _tmp_1492;
  reg [32-1:0] _tmp_1493;
  reg [32-1:0] _tmp_1494;
  reg [32-1:0] _tmp_1495;
  reg [32-1:0] _tmp_1496;
  reg [32-1:0] _tmp_1497;
  reg [32-1:0] _tmp_1498;
  reg [32-1:0] _tmp_1499;
  reg [32-1:0] _tmp_1500;
  reg [32-1:0] _tmp_1501;
  reg [32-1:0] _tmp_1502;
  reg [32-1:0] _tmp_1503;
  reg [32-1:0] _tmp_1504;
  wire [1-1:0] write_rtl_bank_1505;
  assign write_rtl_bank_1505 = _stream_matmul_11_sink_26_sink_waddr;
  assign ram_w16_l512_id0_0_0_addr = (_stream_matmul_11_stream_oready && _stream_matmul_11_sink_26_sink_wenable && (_stream_matmul_11_sink_26_sink_sel == 5) && (write_rtl_bank_1505 == 0))? _stream_matmul_11_sink_26_sink_waddr >> 1 : 
                                     (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_29_source_ram_renable && (_stream_conv2d_4_source_29_source_sel == 12))? _stream_conv2d_4_source_29_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id0_0_0_wdata = (_stream_matmul_11_stream_oready && _stream_matmul_11_sink_26_sink_wenable && (_stream_matmul_11_sink_26_sink_sel == 5) && (write_rtl_bank_1505 == 0))? _stream_matmul_11_sink_26_sink_wdata : 'hx;
  assign ram_w16_l512_id0_0_0_wenable = (_stream_matmul_11_stream_oready && _stream_matmul_11_sink_26_sink_wenable && (_stream_matmul_11_sink_26_sink_sel == 5) && (write_rtl_bank_1505 == 0))? 1'd1 : 0;
  assign ram_w16_l512_id0_0_0_enable = (_stream_matmul_11_stream_oready && _stream_matmul_11_sink_26_sink_wenable && (_stream_matmul_11_sink_26_sink_sel == 5) && (write_rtl_bank_1505 == 0))? 1'd1 : 
                                       (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_29_source_ram_renable && (_stream_conv2d_4_source_29_source_sel == 12))? 1'd1 : 0;
  assign ram_w16_l512_id0_1_0_addr = (_stream_matmul_11_stream_oready && _stream_matmul_11_sink_26_sink_wenable && (_stream_matmul_11_sink_26_sink_sel == 5) && (write_rtl_bank_1505 == 1))? _stream_matmul_11_sink_26_sink_waddr >> 1 : 
                                     (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_29_source_ram_renable && (_stream_conv2d_4_source_29_source_sel == 12))? _stream_conv2d_4_source_29_source_ram_raddr >> 1 : 'hx;
  assign ram_w16_l512_id0_1_0_wdata = (_stream_matmul_11_stream_oready && _stream_matmul_11_sink_26_sink_wenable && (_stream_matmul_11_sink_26_sink_sel == 5) && (write_rtl_bank_1505 == 1))? _stream_matmul_11_sink_26_sink_wdata : 'hx;
  assign ram_w16_l512_id0_1_0_wenable = (_stream_matmul_11_stream_oready && _stream_matmul_11_sink_26_sink_wenable && (_stream_matmul_11_sink_26_sink_sel == 5) && (write_rtl_bank_1505 == 1))? 1'd1 : 0;
  assign ram_w16_l512_id0_1_0_enable = (_stream_matmul_11_stream_oready && _stream_matmul_11_sink_26_sink_wenable && (_stream_matmul_11_sink_26_sink_sel == 5) && (write_rtl_bank_1505 == 1))? 1'd1 : 
                                       (_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_29_source_ram_renable && (_stream_conv2d_4_source_29_source_sel == 12))? 1'd1 : 0;
  reg [32-1:0] _stream_matmul_11_sink_26_sink_fsm_4;
  localparam _stream_matmul_11_sink_26_sink_fsm_4_init = 0;
  wire _set_flag_1506;
  assign _set_flag_1506 = matmul_11_comp_fsm == 4;
  assign _stream_matmul_11_run_flag = (_set_flag_1506)? 1 : 0;
  reg _tmp_1507;
  reg _tmp_1508;
  reg _tmp_1509;
  assign _add_tree_15_source_stop = _add_tree_15_stream_oready && 1'd0;
  reg _tmp_1510;
  reg _tmp_1511;
  assign _add_tree_15_sink_start = _tmp_1511;
  reg _tmp_1512;
  reg _tmp_1513;
  assign _add_tree_15_sink_stop = _tmp_1513;
  reg _tmp_1514;
  reg _tmp_1515;
  assign _add_tree_15_sink_busy = _tmp_1515;
  reg _tmp_1516;
  assign _add_tree_15_busy = _add_tree_15_source_busy || _add_tree_15_sink_busy || _add_tree_15_busy_reg;
  reg _tmp_1517;
  reg _tmp_1518;
  reg _tmp_1519;
  reg _tmp_1520;
  reg _tmp_1521;
  reg _tmp_1522;
  reg [1-1:0] __variable_wdata_2161;
  assign stream_matmul_11__reduce_reset_data = __variable_wdata_2161;
  reg _tmp_1523;
  reg _tmp_1524;
  reg _tmp_1525;
  reg _tmp_1526;
  assign _stream_matmul_11_source_stop = _stream_matmul_11_stream_oready && (_stream_matmul_11_source_11_idle && _stream_matmul_11_source_13_idle && _stream_matmul_11_source_15_idle && _stream_matmul_11_source_20_idle && _stream_matmul_11_source_21_idle && _stream_matmul_11_source_7_idle && _stream_matmul_11_source_9_idle && (_stream_matmul_11_fsm == 3));
  localparam _tmp_1527 = 1;
  wire [_tmp_1527-1:0] _tmp_1528;
  assign _tmp_1528 = _stream_matmul_11_source_11_idle && _stream_matmul_11_source_13_idle && _stream_matmul_11_source_15_idle && _stream_matmul_11_source_20_idle && _stream_matmul_11_source_21_idle && _stream_matmul_11_source_7_idle && _stream_matmul_11_source_9_idle && (_stream_matmul_11_fsm == 3);
  reg [_tmp_1527-1:0] _tmp_1529;
  localparam _tmp_1530 = 1;
  wire [_tmp_1530-1:0] _tmp_1531;
  assign _tmp_1531 = _stream_matmul_11_source_11_idle && _stream_matmul_11_source_13_idle && _stream_matmul_11_source_15_idle && _stream_matmul_11_source_20_idle && _stream_matmul_11_source_21_idle && _stream_matmul_11_source_7_idle && _stream_matmul_11_source_9_idle && (_stream_matmul_11_fsm == 3);
  reg [_tmp_1530-1:0] _tmp_1532;
  reg _tmp_1533;
  reg _tmp_1534;
  reg _tmp_1535;
  reg _tmp_1536;
  reg _tmp_1537;
  reg _tmp_1538;
  reg _tmp_1539;
  reg _tmp_1540;
  reg _tmp_1541;
  reg _tmp_1542;
  reg _tmp_1543;
  reg _tmp_1544;
  reg _tmp_1545;
  reg _tmp_1546;
  reg _tmp_1547;
  reg _tmp_1548;
  reg _tmp_1549;
  reg _tmp_1550;
  reg _tmp_1551;
  reg _tmp_1552;
  reg _tmp_1553;
  reg _tmp_1554;
  reg _tmp_1555;
  reg _tmp_1556;
  reg _tmp_1557;
  reg _tmp_1558;
  reg _tmp_1559;
  reg _tmp_1560;
  reg _tmp_1561;
  reg _tmp_1562;
  reg _tmp_1563;
  assign _stream_matmul_11_sink_start = _tmp_1563;
  reg _tmp_1564;
  reg _tmp_1565;
  reg _tmp_1566;
  reg _tmp_1567;
  reg _tmp_1568;
  reg _tmp_1569;
  reg _tmp_1570;
  reg _tmp_1571;
  reg _tmp_1572;
  reg _tmp_1573;
  reg _tmp_1574;
  reg _tmp_1575;
  reg _tmp_1576;
  reg _tmp_1577;
  reg _tmp_1578;
  reg _tmp_1579;
  reg _tmp_1580;
  reg _tmp_1581;
  reg _tmp_1582;
  reg _tmp_1583;
  reg _tmp_1584;
  reg _tmp_1585;
  reg _tmp_1586;
  reg _tmp_1587;
  reg _tmp_1588;
  reg _tmp_1589;
  reg _tmp_1590;
  reg _tmp_1591;
  reg _tmp_1592;
  reg _tmp_1593;
  reg _tmp_1594;
  assign _stream_matmul_11_sink_stop = _tmp_1594;
  reg _tmp_1595;
  reg _tmp_1596;
  reg _tmp_1597;
  reg _tmp_1598;
  reg _tmp_1599;
  reg _tmp_1600;
  reg _tmp_1601;
  reg _tmp_1602;
  reg _tmp_1603;
  reg _tmp_1604;
  reg _tmp_1605;
  reg _tmp_1606;
  reg _tmp_1607;
  reg _tmp_1608;
  reg _tmp_1609;
  reg _tmp_1610;
  reg _tmp_1611;
  reg _tmp_1612;
  reg _tmp_1613;
  reg _tmp_1614;
  reg _tmp_1615;
  reg _tmp_1616;
  reg _tmp_1617;
  reg _tmp_1618;
  reg _tmp_1619;
  reg _tmp_1620;
  reg _tmp_1621;
  reg _tmp_1622;
  reg _tmp_1623;
  reg _tmp_1624;
  reg _tmp_1625;
  assign _stream_matmul_11_sink_busy = _tmp_1625;
  reg _tmp_1626;
  assign _stream_matmul_11_busy = _stream_matmul_11_source_busy || _stream_matmul_11_sink_busy || _stream_matmul_11_busy_reg;
  wire matmul_11_dma_out_mask_0;
  assign matmul_11_dma_out_mask_0 = matmul_11_out_row_count + 0 >= cparam_matmul_11_out_num_row;
  wire [32-1:0] _dma_write_packed_high_local_size_1627;
  assign _dma_write_packed_high_local_size_1627 = matmul_11_next_out_write_size >> 1;
  wire [1-1:0] _dma_write_packed_low_local_size_1628;
  assign _dma_write_packed_low_local_size_1628 = matmul_11_next_out_write_size & { 1{ 1'd1 } };
  wire [32-1:0] _dma_write_packed_local_packed_size_1629;
  assign _dma_write_packed_local_packed_size_1629 = (_dma_write_packed_low_local_size_1628 > 0)? _dma_write_packed_high_local_size_1627 + 1 : _dma_write_packed_high_local_size_1627;
  wire [32-1:0] mask_addr_shifted_1630;
  assign mask_addr_shifted_1630 = matmul_11_objaddr + (matmul_11_out_base_offset + cparam_matmul_11_out_offset_values_0) + _maxi_global_base_addr >> 2;
  wire [32-1:0] mask_addr_masked_1631;
  assign mask_addr_masked_1631 = mask_addr_shifted_1630 << 2;
  reg [32-1:0] read_burst_packed_fsm_61;
  localparam read_burst_packed_fsm_61_init = 0;
  reg [9-1:0] read_burst_packed_addr_1632;
  reg [9-1:0] read_burst_packed_stride_1633;
  reg [33-1:0] read_burst_packed_length_1634;
  reg read_burst_packed_rvalid_1635;
  reg read_burst_packed_rlast_1636;
  wire [8-1:0] read_burst_packed_ram_addr_1637;
  assign read_burst_packed_ram_addr_1637 = read_burst_packed_addr_1632 >> 1;
  assign ram_w16_l512_id0_0_1_addr = ((read_burst_packed_fsm_61 == 1) && (!read_burst_packed_rvalid_1635 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? read_burst_packed_ram_addr_1637 : 
                                     ((write_burst_packed_fsm_33 == 1) && write_burst_block_ram_wvalid_108)? write_burst_packed_ram_addr_114 : 'hx;
  assign ram_w16_l512_id0_0_1_enable = ((read_burst_packed_fsm_61 == 1) && (!read_burst_packed_rvalid_1635 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? 1'd1 : 
                                       ((write_burst_packed_fsm_33 == 1) && write_burst_block_ram_wvalid_108)? 1'd1 : 0;
  localparam _tmp_1638 = 1;
  wire [_tmp_1638-1:0] _tmp_1639;
  assign _tmp_1639 = (read_burst_packed_fsm_61 == 1) && (!read_burst_packed_rvalid_1635 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0));
  reg [_tmp_1638-1:0] __tmp_1639_1;
  wire [16-1:0] read_burst_packed_ram_rdata_1640;
  assign read_burst_packed_ram_rdata_1640 = ram_w16_l512_id0_0_1_rdata;
  wire [8-1:0] read_burst_packed_ram_addr_1641;
  assign read_burst_packed_ram_addr_1641 = read_burst_packed_addr_1632 >> 1;
  assign ram_w16_l512_id0_1_1_addr = ((read_burst_packed_fsm_61 == 1) && (!read_burst_packed_rvalid_1635 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? read_burst_packed_ram_addr_1641 : 
                                     ((write_burst_packed_fsm_33 == 1) && write_burst_block_ram_wvalid_108)? write_burst_packed_ram_addr_116 : 'hx;
  assign ram_w16_l512_id0_1_1_enable = ((read_burst_packed_fsm_61 == 1) && (!read_burst_packed_rvalid_1635 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)))? 1'd1 : 
                                       ((write_burst_packed_fsm_33 == 1) && write_burst_block_ram_wvalid_108)? 1'd1 : 0;
  localparam _tmp_1642 = 1;
  wire [_tmp_1642-1:0] _tmp_1643;
  assign _tmp_1643 = (read_burst_packed_fsm_61 == 1) && (!read_burst_packed_rvalid_1635 || (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0));
  reg [_tmp_1642-1:0] __tmp_1643_1;
  wire [16-1:0] read_burst_packed_ram_rdata_1644;
  assign read_burst_packed_ram_rdata_1644 = ram_w16_l512_id0_1_1_rdata;
  wire [32-1:0] read_burst_packed_rdata_1645;
  assign read_burst_packed_rdata_1645 = { read_burst_packed_ram_rdata_1644, read_burst_packed_ram_rdata_1640 };
  assign _maxi_write_req_fifo_deq = ((_maxi_write_data_fsm == 2) && (!_maxi_write_req_fifo_empty && (_maxi_write_size_buf == 0)) && !_maxi_write_req_fifo_empty)? 1 : 
                                    ((_maxi_write_data_fsm == 0) && (!_maxi_write_data_busy && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 3)) && !_maxi_write_req_fifo_empty)? 1 : 
                                    ((_maxi_write_data_fsm == 2) && (!_maxi_write_req_fifo_empty && (_maxi_write_size_buf == 0)) && !_maxi_write_req_fifo_empty)? 1 : 
                                    ((_maxi_write_data_fsm == 0) && (!_maxi_write_data_busy && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 2)) && !_maxi_write_req_fifo_empty)? 1 : 
                                    ((_maxi_write_data_fsm == 2) && (!_maxi_write_req_fifo_empty && (_maxi_write_size_buf == 0)) && !_maxi_write_req_fifo_empty)? 1 : 
                                    ((_maxi_write_data_fsm == 0) && (!_maxi_write_data_busy && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 1)) && !_maxi_write_req_fifo_empty)? 1 : 0;
  reg _maxi_wdata_cond_2_1;
  wire matmul_11_update_filter;
  assign matmul_11_update_filter = (cparam_matmul_11_data_stationary == 0) && (matmul_11_row_count >= cparam_matmul_11_max_row_count) && (matmul_11_bat_count >= cparam_matmul_11_max_bat_count) || (cparam_matmul_11_data_stationary == 1) && !cparam_matmul_11_keep_filter;
  wire matmul_11_update_act;
  assign matmul_11_update_act = (cparam_matmul_11_data_stationary == 1) && (matmul_11_och_count >= cparam_matmul_11_max_och_count) || (cparam_matmul_11_data_stationary == 0);
  wire matmul_11_mux_next_dma_flag_0;
  assign matmul_11_mux_next_dma_flag_0 = (matmul_11_row_select == 0)? (matmul_11_row_count >= cparam_matmul_11_max_row_count)? 1 : cparam_matmul_11_dma_flag_conds_0 : 1'd0;

  always @(posedge CLK) begin
    _RESETN_inv_1 <= RESETN_inv;
    _RESETN_inv_2 <= _RESETN_inv_1;
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      maxi_awaddr <= 0;
      maxi_awlen <= 0;
      maxi_awvalid <= 0;
      _maxi_waddr_cond_0_1 <= 0;
    end else begin
      if(_maxi_waddr_cond_0_1) begin
        maxi_awvalid <= 0;
      end 
      if((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (_maxi_outstanding_wcount < 6) && ((_maxi_outstanding_wcount < 6) && (maxi_awready || !maxi_awvalid))) begin
        maxi_awaddr <= _maxi_write_global_addr;
        maxi_awlen <= _maxi_write_cur_global_size - 1;
        maxi_awvalid <= 1;
      end 
      if((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (_maxi_outstanding_wcount < 6) && ((_maxi_outstanding_wcount < 6) && (maxi_awready || !maxi_awvalid)) && (_maxi_write_cur_global_size == 0)) begin
        maxi_awvalid <= 0;
      end 
      _maxi_waddr_cond_0_1 <= 1;
      if(maxi_awvalid && !maxi_awready) begin
        maxi_awvalid <= maxi_awvalid;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _maxi_wdata_sb_0 <= 0;
      _maxi_wvalid_sb_0 <= 0;
      _maxi_wlast_sb_0 <= 0;
      _maxi_wstrb_sb_0 <= 0;
      _maxi_wdata_cond_0_1 <= 0;
      _maxi_wdata_cond_1_1 <= 0;
      _maxi_wdata_cond_2_1 <= 0;
    end else begin
      if(_maxi_wdata_cond_0_1) begin
        _maxi_wvalid_sb_0 <= 0;
        _maxi_wlast_sb_0 <= 0;
      end 
      if(_maxi_wdata_cond_1_1) begin
        _maxi_wvalid_sb_0 <= 0;
        _maxi_wlast_sb_0 <= 0;
      end 
      if(_maxi_wdata_cond_2_1) begin
        _maxi_wvalid_sb_0 <= 0;
        _maxi_wlast_sb_0 <= 0;
      end 
      if((_maxi_write_op_sel_buf == 1) && read_burst_packed_rvalid_1169 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)) && (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0)) begin
        _maxi_wdata_sb_0 <= read_burst_packed_rdata_1179;
        _maxi_wvalid_sb_0 <= 1;
        _maxi_wlast_sb_0 <= read_burst_packed_rlast_1170 || (_maxi_write_size_buf == 1);
        _maxi_wstrb_sb_0 <= { 4{ 1'd1 } };
      end 
      _maxi_wdata_cond_0_1 <= 1;
      if(_maxi_wvalid_sb_0 && !_maxi_wready_sb_0) begin
        _maxi_wvalid_sb_0 <= _maxi_wvalid_sb_0;
        _maxi_wlast_sb_0 <= _maxi_wlast_sb_0;
      end 
      if((_maxi_write_op_sel_buf == 2) && read_burst_packed_rvalid_1301 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)) && (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0)) begin
        _maxi_wdata_sb_0 <= read_burst_packed_rdata_1311;
        _maxi_wvalid_sb_0 <= 1;
        _maxi_wlast_sb_0 <= read_burst_packed_rlast_1302 || (_maxi_write_size_buf == 1);
        _maxi_wstrb_sb_0 <= { 4{ 1'd1 } };
      end 
      _maxi_wdata_cond_1_1 <= 1;
      if(_maxi_wvalid_sb_0 && !_maxi_wready_sb_0) begin
        _maxi_wvalid_sb_0 <= _maxi_wvalid_sb_0;
        _maxi_wlast_sb_0 <= _maxi_wlast_sb_0;
      end 
      if((_maxi_write_op_sel_buf == 3) && read_burst_packed_rvalid_1635 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)) && (_maxi_wready_sb_0 || !_maxi_wvalid_sb_0)) begin
        _maxi_wdata_sb_0 <= read_burst_packed_rdata_1645;
        _maxi_wvalid_sb_0 <= 1;
        _maxi_wlast_sb_0 <= read_burst_packed_rlast_1636 || (_maxi_write_size_buf == 1);
        _maxi_wstrb_sb_0 <= { 4{ 1'd1 } };
      end 
      _maxi_wdata_cond_2_1 <= 1;
      if(_maxi_wvalid_sb_0 && !_maxi_wready_sb_0) begin
        _maxi_wvalid_sb_0 <= _maxi_wvalid_sb_0;
        _maxi_wlast_sb_0 <= _maxi_wlast_sb_0;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _sb_maxi_writedata_data_6 <= 0;
      _sb_maxi_writedata_valid_7 <= 0;
      _sb_maxi_writedata_tmp_data_9 <= 0;
      _sb_maxi_writedata_tmp_valid_10 <= 0;
    end else begin
      if(_sb_maxi_writedata_m_ready_5 || !_sb_maxi_writedata_valid_7) begin
        _sb_maxi_writedata_data_6 <= _sb_maxi_writedata_next_data_11;
        _sb_maxi_writedata_valid_7 <= _sb_maxi_writedata_next_valid_12;
      end 
      if(!_sb_maxi_writedata_tmp_valid_10 && _sb_maxi_writedata_valid_7 && !_sb_maxi_writedata_m_ready_5) begin
        _sb_maxi_writedata_tmp_data_9 <= _sb_maxi_writedata_s_data_3;
        _sb_maxi_writedata_tmp_valid_10 <= _sb_maxi_writedata_s_valid_4;
      end 
      if(_sb_maxi_writedata_tmp_valid_10 && _sb_maxi_writedata_m_ready_5) begin
        _sb_maxi_writedata_tmp_valid_10 <= 0;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      maxi_araddr <= 0;
      maxi_arlen <= 0;
      maxi_arvalid <= 0;
      _maxi_raddr_cond_0_1 <= 0;
    end else begin
      if(_maxi_raddr_cond_0_1) begin
        maxi_arvalid <= 0;
      end 
      if((_maxi_read_req_fsm == 1) && (maxi_arready || !maxi_arvalid)) begin
        maxi_araddr <= _maxi_read_global_addr;
        maxi_arlen <= _maxi_read_cur_global_size - 1;
        maxi_arvalid <= 1;
      end 
      _maxi_raddr_cond_0_1 <= 1;
      if(maxi_arvalid && !maxi_arready) begin
        maxi_arvalid <= maxi_arvalid;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _sb_maxi_readdata_data_21 <= 0;
      _sb_maxi_readdata_valid_22 <= 0;
      _sb_maxi_readdata_tmp_data_24 <= 0;
      _sb_maxi_readdata_tmp_valid_25 <= 0;
    end else begin
      if(_sb_maxi_readdata_m_ready_20 || !_sb_maxi_readdata_valid_22) begin
        _sb_maxi_readdata_data_21 <= _sb_maxi_readdata_next_data_26;
        _sb_maxi_readdata_valid_22 <= _sb_maxi_readdata_next_valid_27;
      end 
      if(!_sb_maxi_readdata_tmp_valid_25 && _sb_maxi_readdata_valid_22 && !_sb_maxi_readdata_m_ready_20) begin
        _sb_maxi_readdata_tmp_data_24 <= _sb_maxi_readdata_s_data_18;
        _sb_maxi_readdata_tmp_valid_25 <= _sb_maxi_readdata_s_valid_19;
      end 
      if(_sb_maxi_readdata_tmp_valid_25 && _sb_maxi_readdata_m_ready_20) begin
        _sb_maxi_readdata_tmp_valid_25 <= 0;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _maxi_outstanding_wcount <= 0;
      _maxi_read_start <= 0;
      _maxi_write_start <= 0;
      _maxi_global_base_addr <= 0;
      _maxi_read_op_sel <= 0;
      _maxi_read_global_addr <= 0;
      _maxi_read_global_size <= 0;
      _maxi_read_local_addr <= 0;
      _maxi_read_local_stride <= 0;
      _maxi_read_local_size <= 0;
      _maxi_read_local_blocksize <= 0;
      _maxi_read_req_busy <= 0;
      _maxi_read_cur_global_size <= 0;
      _maxi_read_data_busy <= 0;
      _maxi_read_op_sel_buf <= 0;
      _maxi_read_local_addr_buf <= 0;
      _maxi_read_local_stride_buf <= 0;
      _maxi_read_local_size_buf <= 0;
      _maxi_read_local_blocksize_buf <= 0;
      _maxi_write_op_sel <= 0;
      _maxi_write_global_addr <= 0;
      _maxi_write_global_size <= 0;
      _maxi_write_local_addr <= 0;
      _maxi_write_local_stride <= 0;
      _maxi_write_local_size <= 0;
      _maxi_write_local_blocksize <= 0;
      _maxi_write_req_busy <= 0;
      _maxi_write_cur_global_size <= 0;
      _maxi_write_data_busy <= 0;
      _maxi_write_op_sel_buf <= 0;
      _maxi_write_local_addr_buf <= 0;
      _maxi_write_local_stride_buf <= 0;
      _maxi_write_size_buf <= 0;
      _maxi_write_local_blocksize_buf <= 0;
    end else begin
      if(maxi_awvalid && maxi_awready && !(maxi_bvalid && maxi_bready) && (_maxi_outstanding_wcount < 7)) begin
        _maxi_outstanding_wcount <= _maxi_outstanding_wcount + 1;
      end 
      if(!(maxi_awvalid && maxi_awready) && (maxi_bvalid && maxi_bready) && (_maxi_outstanding_wcount > 0)) begin
        _maxi_outstanding_wcount <= _maxi_outstanding_wcount - 1;
      end 
      _maxi_read_start <= 0;
      _maxi_write_start <= 0;
      _maxi_global_base_addr <= _saxi_register_32;
      if((control_conv2d_4 == 2) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 1;
        _maxi_read_global_addr <= mask_addr_masked_58;
        _maxi_read_global_size <= _dma_read_packed_local_packed_size_56;
        _maxi_read_local_addr <= 0;
        _maxi_read_local_stride <= 2;
        _maxi_read_local_size <= _dma_read_packed_local_packed_size_56;
        _maxi_read_local_blocksize <= 1;
      end 
      if((_maxi_read_req_fsm == 0) && _maxi_read_start) begin
        _maxi_read_req_busy <= 1;
      end 
      if(_maxi_read_start && _maxi_read_req_fifo_almost_full) begin
        _maxi_read_start <= 1;
      end 
      if((_maxi_read_req_fsm == 0) && (_maxi_read_start || _maxi_read_cont) && !_maxi_read_req_fifo_almost_full && (_maxi_read_global_size <= 256) && ((mask_addr_masked_68 & 4095) + (_maxi_read_global_size << 2) >= 4096)) begin
        _maxi_read_cur_global_size <= 4096 - (mask_addr_masked_70 & 4095) >> 2;
        _maxi_read_global_size <= _maxi_read_global_size - (4096 - (mask_addr_masked_72 & 4095) >> 2);
      end else if((_maxi_read_req_fsm == 0) && (_maxi_read_start || _maxi_read_cont) && !_maxi_read_req_fifo_almost_full && (_maxi_read_global_size <= 256)) begin
        _maxi_read_cur_global_size <= _maxi_read_global_size;
        _maxi_read_global_size <= 0;
      end else if((_maxi_read_req_fsm == 0) && (_maxi_read_start || _maxi_read_cont) && !_maxi_read_req_fifo_almost_full && ((mask_addr_masked_74 & 4095) + 1024 >= 4096)) begin
        _maxi_read_cur_global_size <= 4096 - (mask_addr_masked_76 & 4095) >> 2;
        _maxi_read_global_size <= _maxi_read_global_size - (4096 - (mask_addr_masked_78 & 4095) >> 2);
      end else if((_maxi_read_req_fsm == 0) && (_maxi_read_start || _maxi_read_cont) && !_maxi_read_req_fifo_almost_full) begin
        _maxi_read_cur_global_size <= 256;
        _maxi_read_global_size <= _maxi_read_global_size - 256;
      end 
      if((_maxi_read_req_fsm == 1) && (maxi_arready || !maxi_arvalid)) begin
        _maxi_read_global_addr <= _maxi_read_global_addr + (_maxi_read_cur_global_size << 2);
      end 
      if((_maxi_read_req_fsm == 1) && (maxi_arready || !maxi_arvalid) && (_maxi_read_global_size == 0)) begin
        _maxi_read_req_busy <= 0;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 1))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_conv2d_4 == 4) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 2;
        _maxi_read_global_addr <= mask_addr_masked_91;
        _maxi_read_global_size <= _dma_read_packed_local_packed_size_89;
        _maxi_read_local_addr <= 0;
        _maxi_read_local_stride <= 2;
        _maxi_read_local_size <= _dma_read_packed_local_packed_size_89;
        _maxi_read_local_blocksize <= 1;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 2))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_conv2d_4 == 8) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 3;
        _maxi_read_global_addr <= mask_addr_masked_107;
        _maxi_read_global_size <= _dma_write_block_local_size_102;
        _maxi_read_local_addr <= conv2d_4_filter_page_dma_offset;
        _maxi_read_local_stride <= 2;
        _maxi_read_local_size <= _dma_write_block_local_size_102;
        _maxi_read_local_blocksize <= _dma_read_block_local_blocksize_105;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 3))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_conv2d_4 == 14) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 4;
        _maxi_read_global_addr <= mask_addr_masked_209;
        _maxi_read_global_size <= _dma_write_block_local_size_204;
        _maxi_read_local_addr <= conv2d_4_act_page_dma_offset_0;
        _maxi_read_local_stride <= 2;
        _maxi_read_local_size <= _dma_write_block_local_size_204;
        _maxi_read_local_blocksize <= _dma_read_block_local_blocksize_207;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 4))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_conv2d_4 == 17) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 5;
        _maxi_read_global_addr <= mask_addr_masked_251;
        _maxi_read_global_size <= _dma_write_block_local_size_246;
        _maxi_read_local_addr <= conv2d_4_act_page_dma_offset_1;
        _maxi_read_local_stride <= 2;
        _maxi_read_local_size <= _dma_write_block_local_size_246;
        _maxi_read_local_blocksize <= _dma_read_block_local_blocksize_249;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 5))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_conv2d_4 == 20) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 6;
        _maxi_read_global_addr <= mask_addr_masked_293;
        _maxi_read_global_size <= _dma_write_block_local_size_288;
        _maxi_read_local_addr <= conv2d_4_act_page_dma_offset_2;
        _maxi_read_local_stride <= 2;
        _maxi_read_local_size <= _dma_write_block_local_size_288;
        _maxi_read_local_blocksize <= _dma_read_block_local_blocksize_291;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 6))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_conv2d_4 == 29) && _maxi_write_req_idle) begin
        _maxi_write_start <= 1;
        _maxi_write_op_sel <= 1;
        _maxi_write_global_addr <= mask_addr_masked_1137;
        _maxi_write_global_size <= _dma_write_packed_local_packed_size_1135;
        _maxi_write_local_addr <= conv2d_4_out_laddr_offset + conv2d_4_out_page_dma_offset;
        _maxi_write_local_stride <= 2;
        _maxi_write_local_size <= _dma_write_packed_local_packed_size_1135;
        _maxi_write_local_blocksize <= 1;
      end 
      if((_maxi_write_req_fsm == 0) && _maxi_write_start) begin
        _maxi_write_req_busy <= 1;
      end 
      if(_maxi_write_start && _maxi_write_req_fifo_almost_full) begin
        _maxi_write_start <= 1;
      end 
      if((_maxi_write_req_fsm == 0) && (_maxi_write_start || _maxi_write_cont) && !_maxi_write_req_fifo_almost_full && (_maxi_write_global_size <= 256) && ((mask_addr_masked_1147 & 4095) + (_maxi_write_global_size << 2) >= 4096)) begin
        _maxi_write_cur_global_size <= 4096 - (mask_addr_masked_1149 & 4095) >> 2;
        _maxi_write_global_size <= _maxi_write_global_size - (4096 - (mask_addr_masked_1151 & 4095) >> 2);
      end else if((_maxi_write_req_fsm == 0) && (_maxi_write_start || _maxi_write_cont) && !_maxi_write_req_fifo_almost_full && (_maxi_write_global_size <= 256)) begin
        _maxi_write_cur_global_size <= _maxi_write_global_size;
        _maxi_write_global_size <= 0;
      end else if((_maxi_write_req_fsm == 0) && (_maxi_write_start || _maxi_write_cont) && !_maxi_write_req_fifo_almost_full && ((mask_addr_masked_1153 & 4095) + 1024 >= 4096)) begin
        _maxi_write_cur_global_size <= 4096 - (mask_addr_masked_1155 & 4095) >> 2;
        _maxi_write_global_size <= _maxi_write_global_size - (4096 - (mask_addr_masked_1157 & 4095) >> 2);
      end else if((_maxi_write_req_fsm == 0) && (_maxi_write_start || _maxi_write_cont) && !_maxi_write_req_fifo_almost_full) begin
        _maxi_write_cur_global_size <= 256;
        _maxi_write_global_size <= _maxi_write_global_size - 256;
      end 
      if((_maxi_write_req_fsm == 1) && ((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (maxi_awready || !maxi_awvalid) && (_maxi_outstanding_wcount < 6))) begin
        _maxi_write_global_addr <= _maxi_write_global_addr + (_maxi_write_cur_global_size << 2);
      end 
      if((_maxi_write_req_fsm == 1) && ((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (maxi_awready || !maxi_awvalid) && (_maxi_outstanding_wcount < 6)) && (_maxi_write_global_size == 0)) begin
        _maxi_write_req_busy <= 0;
      end 
      if((_maxi_write_data_fsm == 0) && (!_maxi_write_data_busy && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 1))) begin
        _maxi_write_data_busy <= 1;
        _maxi_write_op_sel_buf <= _maxi_write_op_sel_fifo;
        _maxi_write_local_addr_buf <= _maxi_write_local_addr_fifo;
        _maxi_write_local_stride_buf <= _maxi_write_local_stride_fifo;
        _maxi_write_size_buf <= _maxi_write_size_fifo;
        _maxi_write_local_blocksize_buf <= _maxi_write_local_blocksize_fifo;
      end 
      if(_maxi_write_data_fsm == 1) begin
        _maxi_write_size_buf <= 0;
      end 
      if((_maxi_write_data_fsm == 2) && (!_maxi_write_req_fifo_empty && (_maxi_write_size_buf == 0))) begin
        _maxi_write_size_buf <= _maxi_write_size_fifo;
      end 
      if((_maxi_write_data_fsm == 2) && read_burst_packed_rvalid_1169 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) begin
        _maxi_write_size_buf <= _maxi_write_size_buf - 1;
      end 
      if((_maxi_write_data_fsm == 2) && ((_maxi_write_op_sel_buf == 1) && read_burst_packed_rvalid_1169 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) && read_burst_packed_rlast_1170) begin
        _maxi_write_data_busy <= 0;
      end 
      if((control_max_pool_serial_6 == 5) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 7;
        _maxi_read_global_addr <= mask_addr_masked_1184;
        _maxi_read_global_size <= _dma_read_packed_local_packed_size_1182;
        _maxi_read_local_addr <= max_pool_serial_6_act_page_dma_offset;
        _maxi_read_local_stride <= 2;
        _maxi_read_local_size <= _dma_read_packed_local_packed_size_1182;
        _maxi_read_local_blocksize <= 1;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 7))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_max_pool_serial_6 == 8) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 7;
        _maxi_read_global_addr <= mask_addr_masked_1197;
        _maxi_read_global_size <= _dma_read_packed_local_packed_size_1195;
        _maxi_read_local_addr <= max_pool_serial_6_act_page_dma_offset + cparam_max_pool_serial_6_act_read_size;
        _maxi_read_local_stride <= 2;
        _maxi_read_local_size <= _dma_read_packed_local_packed_size_1195;
        _maxi_read_local_blocksize <= 1;
      end 
      if((control_max_pool_serial_6 == 15) && _maxi_write_req_idle) begin
        _maxi_write_start <= 1;
        _maxi_write_op_sel <= 2;
        _maxi_write_global_addr <= mask_addr_masked_1297;
        _maxi_write_global_size <= _dma_write_packed_local_packed_size_1295;
        _maxi_write_local_addr <= max_pool_serial_6_out_page_dma_offset;
        _maxi_write_local_stride <= 2;
        _maxi_write_local_size <= _dma_write_packed_local_packed_size_1295;
        _maxi_write_local_blocksize <= 1;
      end 
      if((_maxi_write_data_fsm == 0) && (!_maxi_write_data_busy && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 2))) begin
        _maxi_write_data_busy <= 1;
        _maxi_write_op_sel_buf <= _maxi_write_op_sel_fifo;
        _maxi_write_local_addr_buf <= _maxi_write_local_addr_fifo;
        _maxi_write_local_stride_buf <= _maxi_write_local_stride_fifo;
        _maxi_write_size_buf <= _maxi_write_size_fifo;
        _maxi_write_local_blocksize_buf <= _maxi_write_local_blocksize_fifo;
      end 
      if(_maxi_write_data_fsm == 1) begin
        _maxi_write_size_buf <= 0;
      end 
      if((_maxi_write_data_fsm == 2) && (!_maxi_write_req_fifo_empty && (_maxi_write_size_buf == 0))) begin
        _maxi_write_size_buf <= _maxi_write_size_fifo;
      end 
      if((_maxi_write_data_fsm == 2) && read_burst_packed_rvalid_1301 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) begin
        _maxi_write_size_buf <= _maxi_write_size_buf - 1;
      end 
      if((_maxi_write_data_fsm == 2) && ((_maxi_write_op_sel_buf == 2) && read_burst_packed_rvalid_1301 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) && read_burst_packed_rlast_1302) begin
        _maxi_write_data_busy <= 0;
      end 
      if((control_matmul_11 == 2) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 8;
        _maxi_read_global_addr <= mask_addr_masked_1316;
        _maxi_read_global_size <= _dma_read_packed_local_packed_size_1314;
        _maxi_read_local_addr <= 0;
        _maxi_read_local_stride <= 2;
        _maxi_read_local_size <= _dma_read_packed_local_packed_size_1314;
        _maxi_read_local_blocksize <= 1;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 8))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_matmul_11 == 4) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 9;
        _maxi_read_global_addr <= mask_addr_masked_1329;
        _maxi_read_global_size <= _dma_read_packed_local_packed_size_1327;
        _maxi_read_local_addr <= 0;
        _maxi_read_local_stride <= 2;
        _maxi_read_local_size <= _dma_read_packed_local_packed_size_1327;
        _maxi_read_local_blocksize <= 1;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 9))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_matmul_11 == 8) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 7;
        _maxi_read_global_addr <= mask_addr_masked_1342;
        _maxi_read_global_size <= _dma_read_packed_local_packed_size_1340;
        _maxi_read_local_addr <= matmul_11_filter_page_dma_offset;
        _maxi_read_local_stride <= 2;
        _maxi_read_local_size <= _dma_read_packed_local_packed_size_1340;
        _maxi_read_local_blocksize <= 1;
      end 
      if((control_matmul_11 == 14) && _maxi_read_req_idle) begin
        _maxi_read_start <= 1;
        _maxi_read_op_sel <= 10;
        _maxi_read_global_addr <= mask_addr_masked_1347;
        _maxi_read_global_size <= _dma_read_packed_local_packed_size_1345;
        _maxi_read_local_addr <= matmul_11_act_page_dma_offset_0;
        _maxi_read_local_stride <= 2;
        _maxi_read_local_size <= _dma_read_packed_local_packed_size_1345;
        _maxi_read_local_blocksize <= 1;
      end 
      if((_maxi_read_data_fsm == 0) && (!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 10))) begin
        _maxi_read_data_busy <= 1;
        _maxi_read_op_sel_buf <= _maxi_read_op_sel_fifo;
        _maxi_read_local_addr_buf <= _maxi_read_local_addr_fifo;
        _maxi_read_local_stride_buf <= _maxi_read_local_stride_fifo;
        _maxi_read_local_size_buf <= _maxi_read_local_size_fifo;
        _maxi_read_local_blocksize_buf <= _maxi_read_local_blocksize_fifo;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0) begin
        _maxi_read_local_size_buf <= _maxi_read_local_size_buf - 1;
      end 
      if((_maxi_read_data_fsm == 2) && _maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
        _maxi_read_data_busy <= 0;
      end 
      if((control_matmul_11 == 23) && _maxi_write_req_idle) begin
        _maxi_write_start <= 1;
        _maxi_write_op_sel <= 3;
        _maxi_write_global_addr <= mask_addr_masked_1631;
        _maxi_write_global_size <= _dma_write_packed_local_packed_size_1629;
        _maxi_write_local_addr <= matmul_11_out_laddr_offset + matmul_11_out_page_dma_offset;
        _maxi_write_local_stride <= 2;
        _maxi_write_local_size <= _dma_write_packed_local_packed_size_1629;
        _maxi_write_local_blocksize <= 1;
      end 
      if((_maxi_write_data_fsm == 0) && (!_maxi_write_data_busy && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 3))) begin
        _maxi_write_data_busy <= 1;
        _maxi_write_op_sel_buf <= _maxi_write_op_sel_fifo;
        _maxi_write_local_addr_buf <= _maxi_write_local_addr_fifo;
        _maxi_write_local_stride_buf <= _maxi_write_local_stride_fifo;
        _maxi_write_size_buf <= _maxi_write_size_fifo;
        _maxi_write_local_blocksize_buf <= _maxi_write_local_blocksize_fifo;
      end 
      if(_maxi_write_data_fsm == 1) begin
        _maxi_write_size_buf <= 0;
      end 
      if((_maxi_write_data_fsm == 2) && (!_maxi_write_req_fifo_empty && (_maxi_write_size_buf == 0))) begin
        _maxi_write_size_buf <= _maxi_write_size_fifo;
      end 
      if((_maxi_write_data_fsm == 2) && read_burst_packed_rvalid_1635 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) begin
        _maxi_write_size_buf <= _maxi_write_size_buf - 1;
      end 
      if((_maxi_write_data_fsm == 2) && ((_maxi_write_op_sel_buf == 3) && read_burst_packed_rvalid_1635 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) && read_burst_packed_rlast_1636) begin
        _maxi_write_data_busy <= 0;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      count__maxi_read_req_fifo <= 0;
      __tmp_66_1 <= 0;
    end else begin
      if(_maxi_read_req_fifo_enq && !_maxi_read_req_fifo_full && (_maxi_read_req_fifo_deq && !_maxi_read_req_fifo_empty)) begin
        count__maxi_read_req_fifo <= count__maxi_read_req_fifo;
      end else if(_maxi_read_req_fifo_enq && !_maxi_read_req_fifo_full) begin
        count__maxi_read_req_fifo <= count__maxi_read_req_fifo + 1;
      end else if(_maxi_read_req_fifo_deq && !_maxi_read_req_fifo_empty) begin
        count__maxi_read_req_fifo <= count__maxi_read_req_fifo - 1;
      end 
      __tmp_66_1 <= _tmp_66;
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      count__maxi_write_req_fifo <= 0;
      __tmp_1145_1 <= 0;
      __tmp_1165_1 <= 0;
    end else begin
      if(_maxi_write_req_fifo_enq && !_maxi_write_req_fifo_full && (_maxi_write_req_fifo_deq && !_maxi_write_req_fifo_empty)) begin
        count__maxi_write_req_fifo <= count__maxi_write_req_fifo;
      end else if(_maxi_write_req_fifo_enq && !_maxi_write_req_fifo_full) begin
        count__maxi_write_req_fifo <= count__maxi_write_req_fifo + 1;
      end else if(_maxi_write_req_fifo_deq && !_maxi_write_req_fifo_empty) begin
        count__maxi_write_req_fifo <= count__maxi_write_req_fifo - 1;
      end 
      __tmp_1145_1 <= _tmp_1145;
      __tmp_1165_1 <= _tmp_1165;
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      saxi_rdata <= 0;
      saxi_rvalid <= 0;
      _saxi_rdata_cond_0_1 <= 0;
    end else begin
      if(_saxi_rdata_cond_0_1) begin
        saxi_rvalid <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid)) begin
        saxi_rdata <= axislite_rdata_46;
        saxi_rvalid <= 1;
      end 
      _saxi_rdata_cond_0_1 <= 1;
      if(saxi_rvalid && !saxi_rready) begin
        saxi_rvalid <= saxi_rvalid;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      saxi_bvalid <= 0;
      prev_awvalid_43 <= 0;
      prev_arvalid_44 <= 0;
      writevalid_41 <= 0;
      readvalid_42 <= 0;
      addr_40 <= 0;
      _saxi_register_0 <= 0;
      _saxi_flag_0 <= 0;
      _saxi_register_1 <= 0;
      _saxi_flag_1 <= 0;
      _saxi_register_2 <= 0;
      _saxi_flag_2 <= 0;
      _saxi_register_3 <= 0;
      _saxi_flag_3 <= 0;
      _saxi_register_4 <= 0;
      _saxi_flag_4 <= 0;
      _saxi_register_5 <= 0;
      _saxi_flag_5 <= 0;
      _saxi_register_6 <= 0;
      _saxi_flag_6 <= 0;
      _saxi_register_7 <= 0;
      _saxi_flag_7 <= 0;
      _saxi_register_8 <= 0;
      _saxi_flag_8 <= 0;
      _saxi_register_9 <= 0;
      _saxi_flag_9 <= 0;
      _saxi_register_10 <= 0;
      _saxi_flag_10 <= 0;
      _saxi_register_11 <= 0;
      _saxi_flag_11 <= 0;
      _saxi_register_12 <= 0;
      _saxi_flag_12 <= 0;
      _saxi_register_13 <= 0;
      _saxi_flag_13 <= 0;
      _saxi_register_14 <= 0;
      _saxi_flag_14 <= 0;
      _saxi_register_15 <= 0;
      _saxi_flag_15 <= 0;
      _saxi_register_16 <= 0;
      _saxi_flag_16 <= 0;
      _saxi_register_17 <= 0;
      _saxi_flag_17 <= 0;
      _saxi_register_18 <= 0;
      _saxi_flag_18 <= 0;
      _saxi_register_19 <= 0;
      _saxi_flag_19 <= 0;
      _saxi_register_20 <= 0;
      _saxi_flag_20 <= 0;
      _saxi_register_21 <= 0;
      _saxi_flag_21 <= 0;
      _saxi_register_22 <= 0;
      _saxi_flag_22 <= 0;
      _saxi_register_23 <= 0;
      _saxi_flag_23 <= 0;
      _saxi_register_24 <= 0;
      _saxi_flag_24 <= 0;
      _saxi_register_25 <= 0;
      _saxi_flag_25 <= 0;
      _saxi_register_26 <= 0;
      _saxi_flag_26 <= 0;
      _saxi_register_27 <= 0;
      _saxi_flag_27 <= 0;
      _saxi_register_28 <= 0;
      _saxi_flag_28 <= 0;
      _saxi_register_29 <= 0;
      _saxi_flag_29 <= 0;
      _saxi_register_30 <= 0;
      _saxi_flag_30 <= 0;
      _saxi_register_31 <= 1;
      _saxi_flag_31 <= 0;
      _saxi_register_32 <= 0;
      _saxi_flag_32 <= 0;
      _saxi_register_33 <= 0;
      _saxi_flag_33 <= 0;
      _saxi_register_34 <= 0;
      _saxi_flag_34 <= 0;
      _saxi_register_35 <= 0;
      _saxi_flag_35 <= 0;
      _saxi_register_36 <= 0;
      _saxi_flag_36 <= 0;
      _saxi_register_11[0] <= (0 >> 0) & 1'd1;
      _saxi_register_9[0] <= (0 >> 0) & 1'd1;
      _saxi_register_11[1] <= (0 >> 1) & 1'd1;
      _saxi_register_9[1] <= (0 >> 1) & 1'd1;
      _saxi_register_11[2] <= (0 >> 2) & 1'd1;
      _saxi_register_9[2] <= (0 >> 2) & 1'd1;
      _saxi_register_11[3] <= (0 >> 3) & 1'd1;
      _saxi_register_9[3] <= (0 >> 3) & 1'd1;
      _saxi_register_11[4] <= (0 >> 4) & 1'd1;
      _saxi_register_9[4] <= (0 >> 4) & 1'd1;
      _saxi_register_11[5] <= (0 >> 5) & 1'd1;
      _saxi_register_9[5] <= (0 >> 5) & 1'd1;
      _saxi_register_11[6] <= (0 >> 6) & 1'd1;
      _saxi_register_9[6] <= (0 >> 6) & 1'd1;
      _saxi_register_11[7] <= (0 >> 7) & 1'd1;
      _saxi_register_9[7] <= (0 >> 7) & 1'd1;
      _saxi_register_11[8] <= (0 >> 8) & 1'd1;
      _saxi_register_9[8] <= (0 >> 8) & 1'd1;
      _saxi_register_11[9] <= (0 >> 9) & 1'd1;
      _saxi_register_9[9] <= (0 >> 9) & 1'd1;
      _saxi_register_11[10] <= (0 >> 10) & 1'd1;
      _saxi_register_9[10] <= (0 >> 10) & 1'd1;
      _saxi_register_11[11] <= (0 >> 11) & 1'd1;
      _saxi_register_9[11] <= (0 >> 11) & 1'd1;
      _saxi_register_11[12] <= (0 >> 12) & 1'd1;
      _saxi_register_9[12] <= (0 >> 12) & 1'd1;
      _saxi_register_11[13] <= (0 >> 13) & 1'd1;
      _saxi_register_9[13] <= (0 >> 13) & 1'd1;
      _saxi_register_11[14] <= (0 >> 14) & 1'd1;
      _saxi_register_9[14] <= (0 >> 14) & 1'd1;
      _saxi_register_11[15] <= (0 >> 15) & 1'd1;
      _saxi_register_9[15] <= (0 >> 15) & 1'd1;
      _saxi_register_11[16] <= (0 >> 16) & 1'd1;
      _saxi_register_9[16] <= (0 >> 16) & 1'd1;
      _saxi_register_11[17] <= (0 >> 17) & 1'd1;
      _saxi_register_9[17] <= (0 >> 17) & 1'd1;
      _saxi_register_11[18] <= (0 >> 18) & 1'd1;
      _saxi_register_9[18] <= (0 >> 18) & 1'd1;
      _saxi_register_11[19] <= (0 >> 19) & 1'd1;
      _saxi_register_9[19] <= (0 >> 19) & 1'd1;
      _saxi_register_11[20] <= (0 >> 20) & 1'd1;
      _saxi_register_9[20] <= (0 >> 20) & 1'd1;
      _saxi_register_11[21] <= (0 >> 21) & 1'd1;
      _saxi_register_9[21] <= (0 >> 21) & 1'd1;
      _saxi_register_11[22] <= (0 >> 22) & 1'd1;
      _saxi_register_9[22] <= (0 >> 22) & 1'd1;
      _saxi_register_11[23] <= (0 >> 23) & 1'd1;
      _saxi_register_9[23] <= (0 >> 23) & 1'd1;
      _saxi_register_11[24] <= (0 >> 24) & 1'd1;
      _saxi_register_9[24] <= (0 >> 24) & 1'd1;
      _saxi_register_11[25] <= (0 >> 25) & 1'd1;
      _saxi_register_9[25] <= (0 >> 25) & 1'd1;
      _saxi_register_11[26] <= (0 >> 26) & 1'd1;
      _saxi_register_9[26] <= (0 >> 26) & 1'd1;
      _saxi_register_11[27] <= (0 >> 27) & 1'd1;
      _saxi_register_9[27] <= (0 >> 27) & 1'd1;
      _saxi_register_11[28] <= (0 >> 28) & 1'd1;
      _saxi_register_9[28] <= (0 >> 28) & 1'd1;
      _saxi_register_11[29] <= (0 >> 29) & 1'd1;
      _saxi_register_9[29] <= (0 >> 29) & 1'd1;
      _saxi_register_11[30] <= (0 >> 30) & 1'd1;
      _saxi_register_9[30] <= (0 >> 30) & 1'd1;
      _saxi_register_11[31] <= (0 >> 31) & 1'd1;
      _saxi_register_9[31] <= (0 >> 31) & 1'd1;
      internal_state_counter <= 0;
    end else begin
      if(saxi_bvalid && saxi_bready) begin
        saxi_bvalid <= 0;
      end 
      if(saxi_wvalid && saxi_wready) begin
        saxi_bvalid <= 1;
      end 
      prev_awvalid_43 <= saxi_awvalid;
      prev_arvalid_44 <= saxi_arvalid;
      writevalid_41 <= 0;
      readvalid_42 <= 0;
      if(saxi_awready && saxi_awvalid && !saxi_bvalid) begin
        addr_40 <= saxi_awaddr;
        writevalid_41 <= 1;
      end else if(saxi_arready && saxi_arvalid) begin
        addr_40 <= saxi_araddr;
        readvalid_42 <= 1;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 0)) begin
        _saxi_register_0 <= axislite_resetval_48;
        _saxi_flag_0 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 1)) begin
        _saxi_register_1 <= axislite_resetval_48;
        _saxi_flag_1 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 2)) begin
        _saxi_register_2 <= axislite_resetval_48;
        _saxi_flag_2 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 3)) begin
        _saxi_register_3 <= axislite_resetval_48;
        _saxi_flag_3 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 4)) begin
        _saxi_register_4 <= axislite_resetval_48;
        _saxi_flag_4 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 5)) begin
        _saxi_register_5 <= axislite_resetval_48;
        _saxi_flag_5 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 6)) begin
        _saxi_register_6 <= axislite_resetval_48;
        _saxi_flag_6 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 7)) begin
        _saxi_register_7 <= axislite_resetval_48;
        _saxi_flag_7 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 8)) begin
        _saxi_register_8 <= axislite_resetval_48;
        _saxi_flag_8 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 9)) begin
        _saxi_register_9 <= axislite_resetval_48;
        _saxi_flag_9 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 10)) begin
        _saxi_register_10 <= axislite_resetval_48;
        _saxi_flag_10 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 11)) begin
        _saxi_register_11 <= axislite_resetval_48;
        _saxi_flag_11 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 12)) begin
        _saxi_register_12 <= axislite_resetval_48;
        _saxi_flag_12 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 13)) begin
        _saxi_register_13 <= axislite_resetval_48;
        _saxi_flag_13 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 14)) begin
        _saxi_register_14 <= axislite_resetval_48;
        _saxi_flag_14 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 15)) begin
        _saxi_register_15 <= axislite_resetval_48;
        _saxi_flag_15 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 16)) begin
        _saxi_register_16 <= axislite_resetval_48;
        _saxi_flag_16 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 17)) begin
        _saxi_register_17 <= axislite_resetval_48;
        _saxi_flag_17 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 18)) begin
        _saxi_register_18 <= axislite_resetval_48;
        _saxi_flag_18 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 19)) begin
        _saxi_register_19 <= axislite_resetval_48;
        _saxi_flag_19 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 20)) begin
        _saxi_register_20 <= axislite_resetval_48;
        _saxi_flag_20 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 21)) begin
        _saxi_register_21 <= axislite_resetval_48;
        _saxi_flag_21 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 22)) begin
        _saxi_register_22 <= axislite_resetval_48;
        _saxi_flag_22 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 23)) begin
        _saxi_register_23 <= axislite_resetval_48;
        _saxi_flag_23 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 24)) begin
        _saxi_register_24 <= axislite_resetval_48;
        _saxi_flag_24 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 25)) begin
        _saxi_register_25 <= axislite_resetval_48;
        _saxi_flag_25 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 26)) begin
        _saxi_register_26 <= axislite_resetval_48;
        _saxi_flag_26 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 27)) begin
        _saxi_register_27 <= axislite_resetval_48;
        _saxi_flag_27 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 28)) begin
        _saxi_register_28 <= axislite_resetval_48;
        _saxi_flag_28 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 29)) begin
        _saxi_register_29 <= axislite_resetval_48;
        _saxi_flag_29 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 30)) begin
        _saxi_register_30 <= axislite_resetval_48;
        _saxi_flag_30 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 31)) begin
        _saxi_register_31 <= axislite_resetval_48;
        _saxi_flag_31 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 32)) begin
        _saxi_register_32 <= axislite_resetval_48;
        _saxi_flag_32 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 33)) begin
        _saxi_register_33 <= axislite_resetval_48;
        _saxi_flag_33 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 34)) begin
        _saxi_register_34 <= axislite_resetval_48;
        _saxi_flag_34 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 35)) begin
        _saxi_register_35 <= axislite_resetval_48;
        _saxi_flag_35 <= 0;
      end 
      if((_saxi_register_fsm == 1) && (saxi_rready || !saxi_rvalid) && axislite_flag_47 && (axis_maskaddr_45 == 36)) begin
        _saxi_register_36 <= axislite_resetval_48;
        _saxi_flag_36 <= 0;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 0)) begin
        _saxi_register_0 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 1)) begin
        _saxi_register_1 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 2)) begin
        _saxi_register_2 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 3)) begin
        _saxi_register_3 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 4)) begin
        _saxi_register_4 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 5)) begin
        _saxi_register_5 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 6)) begin
        _saxi_register_6 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 7)) begin
        _saxi_register_7 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 8)) begin
        _saxi_register_8 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 9)) begin
        _saxi_register_9 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 10)) begin
        _saxi_register_10 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 11)) begin
        _saxi_register_11 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 12)) begin
        _saxi_register_12 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 13)) begin
        _saxi_register_13 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 14)) begin
        _saxi_register_14 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 15)) begin
        _saxi_register_15 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 16)) begin
        _saxi_register_16 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 17)) begin
        _saxi_register_17 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 18)) begin
        _saxi_register_18 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 19)) begin
        _saxi_register_19 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 20)) begin
        _saxi_register_20 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 21)) begin
        _saxi_register_21 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 22)) begin
        _saxi_register_22 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 23)) begin
        _saxi_register_23 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 24)) begin
        _saxi_register_24 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 25)) begin
        _saxi_register_25 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 26)) begin
        _saxi_register_26 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 27)) begin
        _saxi_register_27 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 28)) begin
        _saxi_register_28 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 29)) begin
        _saxi_register_29 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 30)) begin
        _saxi_register_30 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 31)) begin
        _saxi_register_31 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 32)) begin
        _saxi_register_32 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 33)) begin
        _saxi_register_33 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 34)) begin
        _saxi_register_34 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 35)) begin
        _saxi_register_35 <= saxi_wdata;
      end 
      if((_saxi_register_fsm == 3) && saxi_wvalid && (axis_maskaddr_45 == 36)) begin
        _saxi_register_36 <= saxi_wdata;
      end 
      if(_saxi_register_11[0] == 1) begin
        _saxi_register_11[0] <= 0;
        _saxi_register_9[0] <= 0;
      end 
      if(_saxi_register_11[1] == 1) begin
        _saxi_register_11[1] <= 0;
        _saxi_register_9[1] <= 0;
      end 
      if(_saxi_register_11[2] == 1) begin
        _saxi_register_11[2] <= 0;
        _saxi_register_9[2] <= 0;
      end 
      if(_saxi_register_11[3] == 1) begin
        _saxi_register_11[3] <= 0;
        _saxi_register_9[3] <= 0;
      end 
      if(_saxi_register_11[4] == 1) begin
        _saxi_register_11[4] <= 0;
        _saxi_register_9[4] <= 0;
      end 
      if(_saxi_register_11[5] == 1) begin
        _saxi_register_11[5] <= 0;
        _saxi_register_9[5] <= 0;
      end 
      if(_saxi_register_11[6] == 1) begin
        _saxi_register_11[6] <= 0;
        _saxi_register_9[6] <= 0;
      end 
      if(_saxi_register_11[7] == 1) begin
        _saxi_register_11[7] <= 0;
        _saxi_register_9[7] <= 0;
      end 
      if(_saxi_register_11[8] == 1) begin
        _saxi_register_11[8] <= 0;
        _saxi_register_9[8] <= 0;
      end 
      if(_saxi_register_11[9] == 1) begin
        _saxi_register_11[9] <= 0;
        _saxi_register_9[9] <= 0;
      end 
      if(_saxi_register_11[10] == 1) begin
        _saxi_register_11[10] <= 0;
        _saxi_register_9[10] <= 0;
      end 
      if(_saxi_register_11[11] == 1) begin
        _saxi_register_11[11] <= 0;
        _saxi_register_9[11] <= 0;
      end 
      if(_saxi_register_11[12] == 1) begin
        _saxi_register_11[12] <= 0;
        _saxi_register_9[12] <= 0;
      end 
      if(_saxi_register_11[13] == 1) begin
        _saxi_register_11[13] <= 0;
        _saxi_register_9[13] <= 0;
      end 
      if(_saxi_register_11[14] == 1) begin
        _saxi_register_11[14] <= 0;
        _saxi_register_9[14] <= 0;
      end 
      if(_saxi_register_11[15] == 1) begin
        _saxi_register_11[15] <= 0;
        _saxi_register_9[15] <= 0;
      end 
      if(_saxi_register_11[16] == 1) begin
        _saxi_register_11[16] <= 0;
        _saxi_register_9[16] <= 0;
      end 
      if(_saxi_register_11[17] == 1) begin
        _saxi_register_11[17] <= 0;
        _saxi_register_9[17] <= 0;
      end 
      if(_saxi_register_11[18] == 1) begin
        _saxi_register_11[18] <= 0;
        _saxi_register_9[18] <= 0;
      end 
      if(_saxi_register_11[19] == 1) begin
        _saxi_register_11[19] <= 0;
        _saxi_register_9[19] <= 0;
      end 
      if(_saxi_register_11[20] == 1) begin
        _saxi_register_11[20] <= 0;
        _saxi_register_9[20] <= 0;
      end 
      if(_saxi_register_11[21] == 1) begin
        _saxi_register_11[21] <= 0;
        _saxi_register_9[21] <= 0;
      end 
      if(_saxi_register_11[22] == 1) begin
        _saxi_register_11[22] <= 0;
        _saxi_register_9[22] <= 0;
      end 
      if(_saxi_register_11[23] == 1) begin
        _saxi_register_11[23] <= 0;
        _saxi_register_9[23] <= 0;
      end 
      if(_saxi_register_11[24] == 1) begin
        _saxi_register_11[24] <= 0;
        _saxi_register_9[24] <= 0;
      end 
      if(_saxi_register_11[25] == 1) begin
        _saxi_register_11[25] <= 0;
        _saxi_register_9[25] <= 0;
      end 
      if(_saxi_register_11[26] == 1) begin
        _saxi_register_11[26] <= 0;
        _saxi_register_9[26] <= 0;
      end 
      if(_saxi_register_11[27] == 1) begin
        _saxi_register_11[27] <= 0;
        _saxi_register_9[27] <= 0;
      end 
      if(_saxi_register_11[28] == 1) begin
        _saxi_register_11[28] <= 0;
        _saxi_register_9[28] <= 0;
      end 
      if(_saxi_register_11[29] == 1) begin
        _saxi_register_11[29] <= 0;
        _saxi_register_9[29] <= 0;
      end 
      if(_saxi_register_11[30] == 1) begin
        _saxi_register_11[30] <= 0;
        _saxi_register_9[30] <= 0;
      end 
      if(_saxi_register_11[31] == 1) begin
        _saxi_register_11[31] <= 0;
        _saxi_register_9[31] <= 0;
      end 
      if(irq_busy_edge_51) begin
        _saxi_register_9[0] <= irq_busy_edge_51;
      end 
      if(irq_extern_edge_53) begin
        _saxi_register_9[1] <= irq_extern_edge_53;
      end 
      if(main_fsm == 0) begin
        _saxi_register_5 <= 0;
        _saxi_register_6 <= 0;
        _saxi_register_7 <= 0;
      end 
      if(main_fsm == 1) begin
        internal_state_counter <= 0;
        _saxi_register_12 <= 0;
      end else if(main_fsm == _saxi_register_13) begin
        if(internal_state_counter == _saxi_register_14) begin
          internal_state_counter <= 0;
          _saxi_register_12 <= _saxi_register_12 + 1;
        end else begin
          internal_state_counter <= internal_state_counter + 1;
        end
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_0 <= 1;
        _saxi_flag_0 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_1 <= 1;
        _saxi_flag_1 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_2 <= 1;
        _saxi_flag_2 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_3 <= 1;
        _saxi_flag_3 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_4 <= 1;
        _saxi_flag_4 <= 0;
      end 
      if((main_fsm == 1) && 1) begin
        _saxi_register_5 <= 1;
        _saxi_flag_5 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_6 <= 1;
        _saxi_flag_6 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_7 <= 1;
        _saxi_flag_7 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_8 <= 1;
        _saxi_flag_8 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_9 <= 1;
        _saxi_flag_9 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_10 <= 1;
        _saxi_flag_10 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_11 <= 1;
        _saxi_flag_11 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_12 <= 1;
        _saxi_flag_12 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_13 <= 1;
        _saxi_flag_13 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_14 <= 1;
        _saxi_flag_14 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_15 <= 1;
        _saxi_flag_15 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_16 <= 1;
        _saxi_flag_16 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_17 <= 1;
        _saxi_flag_17 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_18 <= 1;
        _saxi_flag_18 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_19 <= 1;
        _saxi_flag_19 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_20 <= 1;
        _saxi_flag_20 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_21 <= 1;
        _saxi_flag_21 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_22 <= 1;
        _saxi_flag_22 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_23 <= 1;
        _saxi_flag_23 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_24 <= 1;
        _saxi_flag_24 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_25 <= 1;
        _saxi_flag_25 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_26 <= 1;
        _saxi_flag_26 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_27 <= 1;
        _saxi_flag_27 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_28 <= 1;
        _saxi_flag_28 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_29 <= 1;
        _saxi_flag_29 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_30 <= 1;
        _saxi_flag_30 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_31 <= 1;
        _saxi_flag_31 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_32 <= 1;
        _saxi_flag_32 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_33 <= 1;
        _saxi_flag_33 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_34 <= 1;
        _saxi_flag_34 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_35 <= 1;
        _saxi_flag_35 <= 0;
      end 
      if((main_fsm == 1) && 0) begin
        _saxi_register_36 <= 1;
        _saxi_flag_36 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_0 <= 0;
        _saxi_flag_0 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_1 <= 0;
        _saxi_flag_1 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_2 <= 0;
        _saxi_flag_2 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_3 <= 0;
        _saxi_flag_3 <= 0;
      end 
      if((main_fsm == 2) && 1) begin
        _saxi_register_4 <= 0;
        _saxi_flag_4 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_5 <= 0;
        _saxi_flag_5 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_6 <= 0;
        _saxi_flag_6 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_7 <= 0;
        _saxi_flag_7 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_8 <= 0;
        _saxi_flag_8 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_9 <= 0;
        _saxi_flag_9 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_10 <= 0;
        _saxi_flag_10 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_11 <= 0;
        _saxi_flag_11 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_12 <= 0;
        _saxi_flag_12 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_13 <= 0;
        _saxi_flag_13 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_14 <= 0;
        _saxi_flag_14 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_15 <= 0;
        _saxi_flag_15 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_16 <= 0;
        _saxi_flag_16 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_17 <= 0;
        _saxi_flag_17 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_18 <= 0;
        _saxi_flag_18 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_19 <= 0;
        _saxi_flag_19 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_20 <= 0;
        _saxi_flag_20 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_21 <= 0;
        _saxi_flag_21 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_22 <= 0;
        _saxi_flag_22 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_23 <= 0;
        _saxi_flag_23 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_24 <= 0;
        _saxi_flag_24 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_25 <= 0;
        _saxi_flag_25 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_26 <= 0;
        _saxi_flag_26 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_27 <= 0;
        _saxi_flag_27 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_28 <= 0;
        _saxi_flag_28 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_29 <= 0;
        _saxi_flag_29 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_30 <= 0;
        _saxi_flag_30 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_31 <= 0;
        _saxi_flag_31 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_32 <= 0;
        _saxi_flag_32 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_33 <= 0;
        _saxi_flag_33 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_34 <= 0;
        _saxi_flag_34 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_35 <= 0;
        _saxi_flag_35 <= 0;
      end 
      if((main_fsm == 2) && 0) begin
        _saxi_register_36 <= 0;
        _saxi_flag_36 <= 0;
      end 
      if((main_fsm == 43) && 0) begin
        _saxi_register_0 <= 0;
        _saxi_flag_0 <= 0;
      end 
      if((main_fsm == 43) && 0) begin
        _saxi_register_1 <= 0;
        _saxi_flag_1 <= 0;
      end 
      if((main_fsm == 43) && 0) begin
        _saxi_register_2 <= 0;
        _saxi_flag_2 <= 0;
      end 
      if((main_fsm == 43) && 0) begin
        _saxi_register_3 <= 0;
        _saxi_flag_3 <= 0;
      end 
      if((main_fsm == 43) && 0) begin
        _saxi_register_4 <= 0;
        _saxi_flag_4 <= 0;
      end 
      if((main_fsm == 43) && 1) begin
        _saxi_register_5 <= 0;
        _saxi_flag_5 <= 0;
      end 
      if((main_fsm == 43) && 0) begin
        _saxi_register_6 <= 0;
        _saxi_flag_6 <= 0;
      end 
      if((main_fsm == 43) && 0) begin
        _saxi_register_7 <= 0;
        _saxi_flag_7 <= 0;
      end 
      if((main_fsm == 43) && 0) begin
        _saxi_register_8 <= 0;
        _saxi_flag_8 <= 0;
      end 
      if((main_fsm == 43) && 0) begin
        _saxi_register_9 <= 0;
        _saxi_flag_9 <= 0;
      end 
      if((main_fsm == 43) && 0) begin
        _saxi_register_10 <= 0;
        _saxi_flag_10 <= 0;
      end 
      if((main_fsm == 43) && 0) begin
        _saxi_register_11 <= 0;
        _saxi_flag_11 <= 0;
      end 
      if((main_fsm == 43) && 0) begin
        _saxi_register_12 <= 0;
        _saxi_flag_12 <= 0;
      end 
      if((main_fsm == 43) && 0) begin
        _saxi_register_13 <= 0;
        _saxi_flag_13 <= 0;
      end 
      if((main_fsm == 43) && 0) begin
        _saxi_register_14 <= 0;
        _saxi_flag_14 <= 0;
      end 
      if((main_fsm == 43) && 0) begin
        _saxi_register_15 <= 0;
        _saxi_flag_15 <= 0;
      end 
      if((main_fsm == 43) && 0) begin
        _saxi_register_16 <= 0;
        _saxi_flag_16 <= 0;
      end 
      if((main_fsm == 43) && 0) begin
        _saxi_register_17 <= 0;
        _saxi_flag_17 <= 0;
      end 
      if((main_fsm == 43) && 0) begin
        _saxi_register_18 <= 0;
        _saxi_flag_18 <= 0;
      end 
      if((main_fsm == 43) && 0) begin
        _saxi_register_19 <= 0;
        _saxi_flag_19 <= 0;
      end 
      if((main_fsm == 43) && 0) begin
        _saxi_register_20 <= 0;
        _saxi_flag_20 <= 0;
      end 
      if((main_fsm == 43) && 0) begin
        _saxi_register_21 <= 0;
        _saxi_flag_21 <= 0;
      end 
      if((main_fsm == 43) && 0) begin
        _saxi_register_22 <= 0;
        _saxi_flag_22 <= 0;
      end 
      if((main_fsm == 43) && 0) begin
        _saxi_register_23 <= 0;
        _saxi_flag_23 <= 0;
      end 
      if((main_fsm == 43) && 0) begin
        _saxi_register_24 <= 0;
        _saxi_flag_24 <= 0;
      end 
      if((main_fsm == 43) && 0) begin
        _saxi_register_25 <= 0;
        _saxi_flag_25 <= 0;
      end 
      if((main_fsm == 43) && 0) begin
        _saxi_register_26 <= 0;
        _saxi_flag_26 <= 0;
      end 
      if((main_fsm == 43) && 0) begin
        _saxi_register_27 <= 0;
        _saxi_flag_27 <= 0;
      end 
      if((main_fsm == 43) && 0) begin
        _saxi_register_28 <= 0;
        _saxi_flag_28 <= 0;
      end 
      if((main_fsm == 43) && 0) begin
        _saxi_register_29 <= 0;
        _saxi_flag_29 <= 0;
      end 
      if((main_fsm == 43) && 0) begin
        _saxi_register_30 <= 0;
        _saxi_flag_30 <= 0;
      end 
      if((main_fsm == 43) && 0) begin
        _saxi_register_31 <= 0;
        _saxi_flag_31 <= 0;
      end 
      if((main_fsm == 43) && 0) begin
        _saxi_register_32 <= 0;
        _saxi_flag_32 <= 0;
      end 
      if((main_fsm == 43) && 0) begin
        _saxi_register_33 <= 0;
        _saxi_flag_33 <= 0;
      end 
      if((main_fsm == 43) && 0) begin
        _saxi_register_34 <= 0;
        _saxi_flag_34 <= 0;
      end 
      if((main_fsm == 43) && 0) begin
        _saxi_register_35 <= 0;
        _saxi_flag_35 <= 0;
      end 
      if((main_fsm == 43) && 0) begin
        _saxi_register_36 <= 0;
        _saxi_flag_36 <= 0;
      end 
    end
  end

  localparam _saxi_register_fsm_1 = 1;
  localparam _saxi_register_fsm_2 = 2;
  localparam _saxi_register_fsm_3 = 3;
  localparam _saxi_register_fsm_4 = 4;

  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _saxi_register_fsm <= _saxi_register_fsm_init;
      axis_maskaddr_45 <= 0;
    end else begin
      case(_saxi_register_fsm)
        _saxi_register_fsm_init: begin
          if(readvalid_42 || writevalid_41) begin
            axis_maskaddr_45 <= (addr_40 >> _saxi_shift) & _saxi_mask;
          end 
          if(readvalid_42) begin
            _saxi_register_fsm <= _saxi_register_fsm_1;
          end 
          if(writevalid_41) begin
            _saxi_register_fsm <= _saxi_register_fsm_3;
          end 
        end
        _saxi_register_fsm_1: begin
          if(saxi_rready || !saxi_rvalid) begin
            _saxi_register_fsm <= _saxi_register_fsm_2;
          end 
        end
        _saxi_register_fsm_2: begin
          if(saxi_rready && saxi_rvalid) begin
            _saxi_register_fsm <= _saxi_register_fsm_init;
          end 
        end
        _saxi_register_fsm_3: begin
          if(saxi_wvalid) begin
            _saxi_register_fsm <= _saxi_register_fsm_4;
          end 
        end
        _saxi_register_fsm_4: begin
          if(saxi_bready && saxi_bvalid) begin
            _saxi_register_fsm <= _saxi_register_fsm_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    _rst_logic_1 <= rst_logic;
    _rst_logic_2 <= _rst_logic_1;
    RST <= rst_logic | _rst_logic_1 | _rst_logic_2;
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      irq <= 0;
    end else begin
      irq <= |irq_49;
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      irq_busy_edge_50 <= 0;
    end else begin
      irq_busy_edge_50 <= irq_busy;
    end
  end


  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      irq_extern_edge_52 <= 0;
    end else begin
      irq_extern_edge_52 <= irq_extern;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1204_1 <= 0;
      __tmp_1404_1 <= 0;
    end else begin
      __tmp_1204_1 <= _tmp_1204;
      __tmp_1404_1 <= _tmp_1404;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1206_1 <= 0;
      __tmp_1406_1 <= 0;
    end else begin
      __tmp_1206_1 <= _tmp_1206;
      __tmp_1406_1 <= _tmp_1406;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1305_1 <= 0;
      __tmp_1395_1 <= 0;
    end else begin
      __tmp_1305_1 <= _tmp_1305;
      __tmp_1395_1 <= _tmp_1395;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1309_1 <= 0;
      __tmp_1397_1 <= 0;
    end else begin
      __tmp_1309_1 <= _tmp_1309;
      __tmp_1397_1 <= _tmp_1397;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_448_1 <= 0;
      __tmp_1639_1 <= 0;
    end else begin
      __tmp_448_1 <= _tmp_448;
      __tmp_1639_1 <= _tmp_1639;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_450_1 <= 0;
      __tmp_1643_1 <= 0;
    end else begin
      __tmp_450_1 <= _tmp_450;
      __tmp_1643_1 <= _tmp_1643;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_457_1 <= 0;
      __tmp_1366_1 <= 0;
    end else begin
      __tmp_457_1 <= _tmp_457;
      __tmp_1366_1 <= _tmp_1366;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_459_1 <= 0;
      __tmp_1368_1 <= 0;
    end else begin
      __tmp_459_1 <= _tmp_459;
      __tmp_1368_1 <= _tmp_1368;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_466_1 <= 0;
      __tmp_1376_1 <= 0;
    end else begin
      __tmp_466_1 <= _tmp_466;
      __tmp_1376_1 <= _tmp_1376;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_468_1 <= 0;
      __tmp_1378_1 <= 0;
    end else begin
      __tmp_468_1 <= _tmp_468;
      __tmp_1378_1 <= _tmp_1378;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_475_1 <= 0;
    end else begin
      __tmp_475_1 <= _tmp_475;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_477_1 <= 0;
    end else begin
      __tmp_477_1 <= _tmp_477;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_484_1 <= 0;
    end else begin
      __tmp_484_1 <= _tmp_484;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_486_1 <= 0;
    end else begin
      __tmp_486_1 <= _tmp_486;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_493_1 <= 0;
    end else begin
      __tmp_493_1 <= _tmp_493;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_495_1 <= 0;
    end else begin
      __tmp_495_1 <= _tmp_495;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_502_1 <= 0;
    end else begin
      __tmp_502_1 <= _tmp_502;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_504_1 <= 0;
    end else begin
      __tmp_504_1 <= _tmp_504;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_511_1 <= 0;
    end else begin
      __tmp_511_1 <= _tmp_511;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_513_1 <= 0;
    end else begin
      __tmp_513_1 <= _tmp_513;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_520_1 <= 0;
    end else begin
      __tmp_520_1 <= _tmp_520;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_522_1 <= 0;
    end else begin
      __tmp_522_1 <= _tmp_522;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_338_1 <= 0;
    end else begin
      __tmp_338_1 <= _tmp_338;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_340_1 <= 0;
    end else begin
      __tmp_340_1 <= _tmp_340;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_348_1 <= 0;
    end else begin
      __tmp_348_1 <= _tmp_348;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_350_1 <= 0;
    end else begin
      __tmp_350_1 <= _tmp_350;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_367_1 <= 0;
    end else begin
      __tmp_367_1 <= _tmp_367;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_369_1 <= 0;
    end else begin
      __tmp_369_1 <= _tmp_369;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_376_1 <= 0;
    end else begin
      __tmp_376_1 <= _tmp_376;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_378_1 <= 0;
    end else begin
      __tmp_378_1 <= _tmp_378;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_385_1 <= 0;
    end else begin
      __tmp_385_1 <= _tmp_385;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_387_1 <= 0;
    end else begin
      __tmp_387_1 <= _tmp_387;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_394_1 <= 0;
    end else begin
      __tmp_394_1 <= _tmp_394;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_396_1 <= 0;
    end else begin
      __tmp_396_1 <= _tmp_396;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_403_1 <= 0;
    end else begin
      __tmp_403_1 <= _tmp_403;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_405_1 <= 0;
    end else begin
      __tmp_405_1 <= _tmp_405;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_412_1 <= 0;
    end else begin
      __tmp_412_1 <= _tmp_412;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_414_1 <= 0;
    end else begin
      __tmp_414_1 <= _tmp_414;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_421_1 <= 0;
    end else begin
      __tmp_421_1 <= _tmp_421;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_423_1 <= 0;
    end else begin
      __tmp_423_1 <= _tmp_423;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_430_1 <= 0;
    end else begin
      __tmp_430_1 <= _tmp_430;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_432_1 <= 0;
    end else begin
      __tmp_432_1 <= _tmp_432;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_439_1 <= 0;
    end else begin
      __tmp_439_1 <= _tmp_439;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_441_1 <= 0;
    end else begin
      __tmp_441_1 <= _tmp_441;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1173_1 <= 0;
    end else begin
      __tmp_1173_1 <= _tmp_1173;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1177_1 <= 0;
    end else begin
      __tmp_1177_1 <= _tmp_1177;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _acc_14_x_source_ram_renable <= 0;
      _acc_14_x_source_fifo_deq <= 0;
      _acc_14_x_idle <= 1;
      _acc_14_rshift_source_ram_renable <= 0;
      _acc_14_rshift_source_fifo_deq <= 0;
      _acc_14_rshift_idle <= 1;
      _acc_14_sum_sink_wenable <= 0;
      _acc_14_sum_sink_fifo_enq <= 0;
      _acc_14_valid_sink_wenable <= 0;
      _acc_14_valid_sink_fifo_enq <= 0;
      __acc_14_stream_ivalid_1 <= 0;
      __acc_14_stream_ivalid_2 <= 0;
      __acc_14_stream_ivalid_3 <= 0;
      __acc_14_stream_ivalid_4 <= 0;
      __acc_14_stream_ivalid_5 <= 0;
      _greaterthan_data_1283 <= 0;
      _minus_data_1285 <= 0;
      _reduceadd_data_1296 <= 1'sd0;
      _reduceadd_count_1296 <= 0;
      _reduceadd_prev_count_max_1296 <= 0;
      _pulse_data_1298 <= 1'sd0;
      _pulse_count_1298 <= 0;
      _pulse_prev_count_max_1298 <= 0;
      __delay_data_2103__variable_1281 <= 0;
      _sll_data_1287 <= 0;
      __delay_data_2100_greaterthan_1283 <= 0;
      __delay_data_2101_reduceadd_1296 <= 0;
      __delay_data_2104__delay_2103__variable_1281 <= 0;
      __delay_data_2107_pulse_1298 <= 0;
      _cond_data_1293 <= 0;
      __delay_data_2102__delay_2101_reduceadd_1296 <= 0;
      __delay_data_2105__delay_2104__delay_2103__variable_1281 <= 0;
      __delay_data_2108__delay_2107_pulse_1298 <= 0;
      _plus_data_1300 <= 0;
      __delay_data_2106__delay_2105__delay_2104____variable_1281 <= 0;
      __delay_data_2109__delay_2108__delay_2107_pulse_1298 <= 0;
      _sra_data_1301 <= 0;
      __delay_data_2110__delay_2109__delay_2108___pulse_1298 <= 0;
      __variable_wdata_1295 <= 0;
      __variable_wdata_1280 <= 0;
      __variable_wdata_1281 <= 0;
      __variable_wdata_1282 <= 0;
      _tmp_951 <= 0;
      _tmp_952 <= 0;
      _tmp_953 <= 0;
      _tmp_954 <= 0;
      _tmp_955 <= 0;
      _tmp_956 <= 0;
      _tmp_957 <= 0;
      _tmp_958 <= 0;
      _tmp_959 <= 0;
      _tmp_960 <= 0;
      _tmp_961 <= 0;
      _tmp_962 <= 0;
      _tmp_963 <= 0;
      _tmp_964 <= 0;
      _tmp_965 <= 0;
      _tmp_966 <= 0;
      _tmp_967 <= 0;
      _tmp_968 <= 0;
      _tmp_969 <= 0;
      _tmp_970 <= 0;
      _tmp_971 <= 0;
      _tmp_972 <= 0;
      _tmp_973 <= 0;
      _tmp_974 <= 0;
      _tmp_975 <= 0;
      _tmp_976 <= 0;
      _tmp_977 <= 0;
      _tmp_978 <= 0;
      _tmp_979 <= 0;
      _tmp_980 <= 0;
      _tmp_981 <= 0;
      _tmp_982 <= 0;
      _acc_14_busy_reg <= 0;
    end else begin
      if(_acc_14_stream_oready) begin
        _acc_14_x_source_ram_renable <= 0;
        _acc_14_x_source_fifo_deq <= 0;
      end 
      _acc_14_x_idle <= _acc_14_x_idle;
      if(_acc_14_stream_oready) begin
        _acc_14_rshift_source_ram_renable <= 0;
        _acc_14_rshift_source_fifo_deq <= 0;
      end 
      _acc_14_rshift_idle <= _acc_14_rshift_idle;
      if(_acc_14_stream_oready) begin
        _acc_14_sum_sink_wenable <= 0;
        _acc_14_sum_sink_fifo_enq <= 0;
      end 
      if(_acc_14_stream_oready) begin
        _acc_14_valid_sink_wenable <= 0;
        _acc_14_valid_sink_fifo_enq <= 0;
      end 
      if(_acc_14_stream_oready) begin
        __acc_14_stream_ivalid_1 <= _acc_14_stream_ivalid;
      end 
      if(_acc_14_stream_oready) begin
        __acc_14_stream_ivalid_2 <= __acc_14_stream_ivalid_1;
      end 
      if(_acc_14_stream_oready) begin
        __acc_14_stream_ivalid_3 <= __acc_14_stream_ivalid_2;
      end 
      if(_acc_14_stream_oready) begin
        __acc_14_stream_ivalid_4 <= __acc_14_stream_ivalid_3;
      end 
      if(_acc_14_stream_oready) begin
        __acc_14_stream_ivalid_5 <= __acc_14_stream_ivalid_4;
      end 
      if(_acc_14_stream_oready) begin
        _greaterthan_data_1283 <= acc_14_rshift_data > 1'sd0;
      end 
      if(_acc_14_stream_oready) begin
        _minus_data_1285 <= acc_14_rshift_data - 2'sd1;
      end 
      if(_acc_14_stream_ivalid && _acc_14_stream_oready && _reduceadd_reset_cond_1296) begin
        _reduceadd_data_1296 <= 1'sd0;
      end 
      if(_acc_14_stream_ivalid && _acc_14_stream_oready) begin
        _reduceadd_count_1296 <= (_reduceadd_current_count_1296 >= acc_14_size_data - 1)? 0 : _reduceadd_current_count_1296 + 1;
      end 
      if(_acc_14_stream_ivalid && _acc_14_stream_oready) begin
        _reduceadd_prev_count_max_1296 <= _reduceadd_current_count_1296 >= acc_14_size_data - 1;
      end 
      if(_acc_14_stream_ivalid && _acc_14_stream_oready) begin
        _reduceadd_data_1296 <= _reduceadd_current_data_1296 + acc_14_x_data;
      end 
      if(_acc_14_stream_ivalid && _acc_14_stream_oready && _pulse_reset_cond_1298) begin
        _pulse_data_1298 <= 1'sd0;
      end 
      if(_acc_14_stream_ivalid && _acc_14_stream_oready) begin
        _pulse_count_1298 <= (_pulse_current_count_1298 >= acc_14_size_data - 1)? 0 : _pulse_current_count_1298 + 1;
      end 
      if(_acc_14_stream_ivalid && _acc_14_stream_oready) begin
        _pulse_prev_count_max_1298 <= _pulse_current_count_1298 >= acc_14_size_data - 1;
      end 
      if(_acc_14_stream_ivalid && _acc_14_stream_oready) begin
        _pulse_data_1298 <= _pulse_current_count_1298 >= acc_14_size_data - 1;
      end 
      if(_acc_14_stream_oready) begin
        __delay_data_2103__variable_1281 <= acc_14_rshift_data;
      end 
      if(_acc_14_stream_oready) begin
        _sll_data_1287 <= 2'sd1 << _minus_data_1285;
      end 
      if(_acc_14_stream_oready) begin
        __delay_data_2100_greaterthan_1283 <= _greaterthan_data_1283;
      end 
      if(_acc_14_stream_oready) begin
        __delay_data_2101_reduceadd_1296 <= _reduceadd_data_1296;
      end 
      if(_acc_14_stream_oready) begin
        __delay_data_2104__delay_2103__variable_1281 <= __delay_data_2103__variable_1281;
      end 
      if(_acc_14_stream_oready) begin
        __delay_data_2107_pulse_1298 <= _pulse_data_1298;
      end 
      if(_acc_14_stream_oready) begin
        _cond_data_1293 <= (__delay_data_2100_greaterthan_1283)? _sll_data_1287 : 1'sd0;
      end 
      if(_acc_14_stream_oready) begin
        __delay_data_2102__delay_2101_reduceadd_1296 <= __delay_data_2101_reduceadd_1296;
      end 
      if(_acc_14_stream_oready) begin
        __delay_data_2105__delay_2104__delay_2103__variable_1281 <= __delay_data_2104__delay_2103__variable_1281;
      end 
      if(_acc_14_stream_oready) begin
        __delay_data_2108__delay_2107_pulse_1298 <= __delay_data_2107_pulse_1298;
      end 
      if(_acc_14_stream_oready) begin
        _plus_data_1300 <= __delay_data_2102__delay_2101_reduceadd_1296 + _cond_data_1293;
      end 
      if(_acc_14_stream_oready) begin
        __delay_data_2106__delay_2105__delay_2104____variable_1281 <= __delay_data_2105__delay_2104__delay_2103__variable_1281;
      end 
      if(_acc_14_stream_oready) begin
        __delay_data_2109__delay_2108__delay_2107_pulse_1298 <= __delay_data_2108__delay_2107_pulse_1298;
      end 
      if(_acc_14_stream_oready) begin
        _sra_data_1301 <= _plus_data_1300 >>> __delay_data_2106__delay_2105__delay_2104____variable_1281;
      end 
      if(_acc_14_stream_oready) begin
        __delay_data_2110__delay_2109__delay_2108___pulse_1298 <= __delay_data_2109__delay_2108__delay_2107_pulse_1298;
      end 
      if(__stream_conv2d_4_stream_ivalid_13 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_1295 <= __delay_data_2297__delay_2296__delay_2295____variable_1553;
      end 
      if(__stream_conv2d_4_stream_ivalid_13 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_1280 <= __substreamoutput_data_2098;
      end 
      if(__stream_conv2d_4_stream_ivalid_13 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_1281 <= __delay_data_2309__delay_2308__delay_2307___plus_2111;
      end 
      if(__stream_conv2d_4_stream_ivalid_13 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_1282 <= __delay_data_2322__delay_2321__delay_2320____variable_1548;
      end 
      if(_acc_14_stream_oready) begin
        _tmp_951 <= _acc_14_source_start;
      end 
      if(_acc_14_stream_oready) begin
        _tmp_952 <= _tmp_951;
      end 
      if(_acc_14_stream_oready) begin
        _tmp_953 <= _tmp_952;
      end 
      if(_acc_14_stream_oready) begin
        _tmp_954 <= _acc_14_source_start;
      end 
      if(_acc_14_stream_oready) begin
        _tmp_955 <= _tmp_954;
      end 
      if(_acc_14_stream_oready) begin
        _tmp_956 <= _tmp_955;
      end 
      if(_acc_14_stream_oready && _tmp_956) begin
        __variable_wdata_1295 <= 1;
      end 
      if(_acc_14_stream_oready) begin
        _tmp_957 <= _acc_14_source_start;
      end 
      if(_acc_14_stream_oready) begin
        _tmp_958 <= _tmp_957;
      end 
      if(_acc_14_stream_oready) begin
        _tmp_959 <= _tmp_958;
      end 
      if(_acc_14_stream_oready) begin
        _tmp_960 <= _tmp_959;
      end 
      if(_acc_14_stream_oready && _tmp_960) begin
        __variable_wdata_1295 <= 0;
      end 
      if(_acc_14_stream_oready && 1'd0) begin
        __variable_wdata_1295 <= 1;
      end 
      if(_acc_14_stream_oready) begin
        _tmp_961 <= _acc_14_source_start;
      end 
      if(_acc_14_stream_oready) begin
        _tmp_962 <= _tmp_961;
      end 
      if(_acc_14_stream_oready) begin
        _tmp_963 <= _tmp_962;
      end 
      if(_acc_14_stream_oready) begin
        _tmp_964 <= _tmp_963;
      end 
      if(_acc_14_stream_oready) begin
        _tmp_965 <= _tmp_964;
      end 
      if(_acc_14_stream_oready) begin
        _tmp_966 <= _tmp_965;
      end 
      if(_acc_14_stream_oready) begin
        _tmp_967 <= _tmp_966;
      end 
      if(_acc_14_stream_oready) begin
        _tmp_968 <= _acc_14_source_stop;
      end 
      if(_acc_14_stream_oready) begin
        _tmp_969 <= _tmp_968;
      end 
      if(_acc_14_stream_oready) begin
        _tmp_970 <= _tmp_969;
      end 
      if(_acc_14_stream_oready) begin
        _tmp_971 <= _tmp_970;
      end 
      if(_acc_14_stream_oready) begin
        _tmp_972 <= _tmp_971;
      end 
      if(_acc_14_stream_oready) begin
        _tmp_973 <= _tmp_972;
      end 
      if(_acc_14_stream_oready) begin
        _tmp_974 <= _tmp_973;
      end 
      if(_acc_14_stream_oready) begin
        _tmp_975 <= _acc_14_source_busy;
      end 
      if(_acc_14_stream_oready) begin
        _tmp_976 <= _tmp_975;
      end 
      if(_acc_14_stream_oready) begin
        _tmp_977 <= _tmp_976;
      end 
      if(_acc_14_stream_oready) begin
        _tmp_978 <= _tmp_977;
      end 
      if(_acc_14_stream_oready) begin
        _tmp_979 <= _tmp_978;
      end 
      if(_acc_14_stream_oready) begin
        _tmp_980 <= _tmp_979;
      end 
      if(_acc_14_stream_oready) begin
        _tmp_981 <= _tmp_980;
      end 
      if(_acc_14_stream_oready) begin
        _tmp_982 <= _acc_14_sink_busy;
      end 
      if(!_acc_14_sink_busy && _tmp_982) begin
        _acc_14_busy_reg <= 0;
      end 
      if(_acc_14_source_busy) begin
        _acc_14_busy_reg <= 1;
      end 
      if(__stream_matmul_11_stream_ivalid_11 && _stream_matmul_11_stream_oready) begin
        __variable_wdata_1295 <= __delay_data_2416__delay_2415__delay_2414____variable_2161;
      end 
      if(__stream_matmul_11_stream_ivalid_11 && _stream_matmul_11_stream_oready) begin
        __variable_wdata_1280 <= __substreamoutput_data_2238;
      end 
      if(__stream_matmul_11_stream_ivalid_11 && _stream_matmul_11_stream_oready) begin
        __variable_wdata_1281 <= __delay_data_2426__delay_2425__delay_2424___plus_2240;
      end 
      if(__stream_matmul_11_stream_ivalid_11 && _stream_matmul_11_stream_oready) begin
        __variable_wdata_1282 <= __delay_data_2437__delay_2436__delay_2435____variable_2156;
      end 
    end
  end

  localparam _acc_14_fsm_1 = 1;
  localparam _acc_14_fsm_2 = 2;
  localparam _acc_14_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _acc_14_fsm <= _acc_14_fsm_init;
      _acc_14_source_start <= 0;
      _acc_14_source_busy <= 0;
      _acc_14_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_13 && _stream_conv2d_4_stream_oready) begin
        _acc_14_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _acc_14_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_acc_14_stream_oready && _tmp_953) begin
        _acc_14_stream_ivalid <= 1;
      end 
      if(_acc_14_stream_oready && 1'd0) begin
        _acc_14_stream_ivalid <= 0;
      end 
      if(__stream_matmul_11_stream_ivalid_11 && _stream_matmul_11_stream_oready) begin
        _acc_14_stream_ivalid <= 1'd1;
      end 
      if(_stream_matmul_11_stream_oready && _stream_matmul_11_busy) begin
        _acc_14_source_busy <= _stream_matmul_11_source_busy;
      end 
      case(_acc_14_fsm)
        _acc_14_fsm_init: begin
          if(_acc_14_run_flag) begin
            _acc_14_source_start <= 1;
          end 
          if(_acc_14_run_flag) begin
            _acc_14_fsm <= _acc_14_fsm_1;
          end 
        end
        _acc_14_fsm_1: begin
          if(_acc_14_source_start && _acc_14_stream_oready) begin
            _acc_14_source_start <= 0;
            _acc_14_source_busy <= 1;
          end 
          if(_acc_14_source_start && _acc_14_stream_oready) begin
            _acc_14_fsm <= _acc_14_fsm_2;
          end 
        end
        _acc_14_fsm_2: begin
          if(_acc_14_stream_oready) begin
            _acc_14_fsm <= _acc_14_fsm_3;
          end 
        end
        _acc_14_fsm_3: begin
          if(_acc_14_stream_oready && 1'd0) begin
            _acc_14_source_busy <= 0;
          end 
          if(_acc_14_stream_oready && 1'd0 && _acc_14_run_flag) begin
            _acc_14_source_start <= 1;
          end 
          if(_acc_14_stream_oready && 1'd0) begin
            _acc_14_fsm <= _acc_14_fsm_init;
          end 
          if(_acc_14_stream_oready && 1'd0 && _acc_14_run_flag) begin
            _acc_14_fsm <= _acc_14_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _add_tree_15_var0_source_ram_renable <= 0;
      _add_tree_15_var0_source_fifo_deq <= 0;
      _add_tree_15_var0_idle <= 1;
      _add_tree_15_sum_sink_wenable <= 0;
      _add_tree_15_sum_sink_fifo_enq <= 0;
      __variable_wdata_1302 <= 0;
      _tmp_1507 <= 0;
      _tmp_1508 <= 0;
      _tmp_1509 <= 0;
      _tmp_1510 <= 0;
      _tmp_1511 <= 0;
      _tmp_1512 <= 0;
      _tmp_1513 <= 0;
      _tmp_1514 <= 0;
      _tmp_1515 <= 0;
      _tmp_1516 <= 0;
      _add_tree_15_busy_reg <= 0;
    end else begin
      if(_add_tree_15_stream_oready) begin
        _add_tree_15_var0_source_ram_renable <= 0;
        _add_tree_15_var0_source_fifo_deq <= 0;
      end 
      _add_tree_15_var0_idle <= _add_tree_15_var0_idle;
      if(_add_tree_15_stream_oready) begin
        _add_tree_15_sum_sink_wenable <= 0;
        _add_tree_15_sum_sink_fifo_enq <= 0;
      end 
      if(__stream_matmul_11_stream_ivalid_10 && _stream_matmul_11_stream_oready) begin
        __variable_wdata_1302 <= __substreamoutput_data_2236;
      end 
      if(_add_tree_15_stream_oready) begin
        _tmp_1507 <= _add_tree_15_source_start;
      end 
      if(_add_tree_15_stream_oready) begin
        _tmp_1508 <= _tmp_1507;
      end 
      if(_add_tree_15_stream_oready) begin
        _tmp_1509 <= _tmp_1508;
      end 
      if(_add_tree_15_stream_oready) begin
        _tmp_1510 <= _add_tree_15_source_start;
      end 
      if(_add_tree_15_stream_oready) begin
        _tmp_1511 <= _tmp_1510;
      end 
      if(_add_tree_15_stream_oready) begin
        _tmp_1512 <= _add_tree_15_source_stop;
      end 
      if(_add_tree_15_stream_oready) begin
        _tmp_1513 <= _tmp_1512;
      end 
      if(_add_tree_15_stream_oready) begin
        _tmp_1514 <= _add_tree_15_source_busy;
      end 
      if(_add_tree_15_stream_oready) begin
        _tmp_1515 <= _tmp_1514;
      end 
      if(_add_tree_15_stream_oready) begin
        _tmp_1516 <= _add_tree_15_sink_busy;
      end 
      if(!_add_tree_15_sink_busy && _tmp_1516) begin
        _add_tree_15_busy_reg <= 0;
      end 
      if(_add_tree_15_source_busy) begin
        _add_tree_15_busy_reg <= 1;
      end 
    end
  end

  localparam _add_tree_15_fsm_1 = 1;
  localparam _add_tree_15_fsm_2 = 2;
  localparam _add_tree_15_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _add_tree_15_fsm <= _add_tree_15_fsm_init;
      _add_tree_15_source_start <= 0;
      _add_tree_15_source_busy <= 0;
      _add_tree_15_stream_ivalid <= 0;
    end else begin
      if(__stream_matmul_11_stream_ivalid_10 && _stream_matmul_11_stream_oready) begin
        _add_tree_15_stream_ivalid <= 1'd1;
      end 
      if(_stream_matmul_11_stream_oready && _stream_matmul_11_busy) begin
        _add_tree_15_source_busy <= _stream_matmul_11_source_busy;
      end 
      if(_add_tree_15_stream_oready && _tmp_1509) begin
        _add_tree_15_stream_ivalid <= 1;
      end 
      if(_add_tree_15_stream_oready && 1'd0) begin
        _add_tree_15_stream_ivalid <= 0;
      end 
      case(_add_tree_15_fsm)
        _add_tree_15_fsm_init: begin
          if(_add_tree_15_run_flag) begin
            _add_tree_15_source_start <= 1;
          end 
          if(_add_tree_15_run_flag) begin
            _add_tree_15_fsm <= _add_tree_15_fsm_1;
          end 
        end
        _add_tree_15_fsm_1: begin
          if(_add_tree_15_source_start && _add_tree_15_stream_oready) begin
            _add_tree_15_source_start <= 0;
            _add_tree_15_source_busy <= 1;
          end 
          if(_add_tree_15_source_start && _add_tree_15_stream_oready) begin
            _add_tree_15_fsm <= _add_tree_15_fsm_2;
          end 
        end
        _add_tree_15_fsm_2: begin
          if(_add_tree_15_stream_oready) begin
            _add_tree_15_fsm <= _add_tree_15_fsm_3;
          end 
        end
        _add_tree_15_fsm_3: begin
          if(_add_tree_15_stream_oready && 1'd0) begin
            _add_tree_15_source_busy <= 0;
          end 
          if(_add_tree_15_stream_oready && 1'd0 && _add_tree_15_run_flag) begin
            _add_tree_15_source_start <= 1;
          end 
          if(_add_tree_15_stream_oready && 1'd0) begin
            _add_tree_15_fsm <= _add_tree_15_fsm_init;
          end 
          if(_add_tree_15_stream_oready && 1'd0 && _add_tree_15_run_flag) begin
            _add_tree_15_fsm <= _add_tree_15_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _add_tree_16_var0_source_ram_renable <= 0;
      _add_tree_16_var0_source_fifo_deq <= 0;
      _add_tree_16_var0_idle <= 1;
      _add_tree_16_var1_source_ram_renable <= 0;
      _add_tree_16_var1_source_fifo_deq <= 0;
      _add_tree_16_var1_idle <= 1;
      _add_tree_16_var2_source_ram_renable <= 0;
      _add_tree_16_var2_source_fifo_deq <= 0;
      _add_tree_16_var2_idle <= 1;
      _add_tree_16_var3_source_ram_renable <= 0;
      _add_tree_16_var3_source_fifo_deq <= 0;
      _add_tree_16_var3_idle <= 1;
      _add_tree_16_var4_source_ram_renable <= 0;
      _add_tree_16_var4_source_fifo_deq <= 0;
      _add_tree_16_var4_idle <= 1;
      _add_tree_16_var5_source_ram_renable <= 0;
      _add_tree_16_var5_source_fifo_deq <= 0;
      _add_tree_16_var5_idle <= 1;
      _add_tree_16_var6_source_ram_renable <= 0;
      _add_tree_16_var6_source_fifo_deq <= 0;
      _add_tree_16_var6_idle <= 1;
      _add_tree_16_var7_source_ram_renable <= 0;
      _add_tree_16_var7_source_fifo_deq <= 0;
      _add_tree_16_var7_idle <= 1;
      _add_tree_16_var8_source_ram_renable <= 0;
      _add_tree_16_var8_source_fifo_deq <= 0;
      _add_tree_16_var8_idle <= 1;
      _add_tree_16_sum_sink_wenable <= 0;
      _add_tree_16_sum_sink_fifo_enq <= 0;
      __add_tree_16_stream_ivalid_1 <= 0;
      __add_tree_16_stream_ivalid_2 <= 0;
      __plusn_data_1314 <= 0;
      __plusn_data_1315 <= 0;
      __plusn_data_1316 <= 0;
      __plusn_data_1317 <= 0;
      __variable_wdata_1304 <= 0;
      __variable_wdata_1305 <= 0;
      __variable_wdata_1306 <= 0;
      __variable_wdata_1307 <= 0;
      __variable_wdata_1308 <= 0;
      __variable_wdata_1309 <= 0;
      __variable_wdata_1310 <= 0;
      __variable_wdata_1311 <= 0;
      __variable_wdata_1312 <= 0;
      _tmp_935 <= 0;
      _tmp_936 <= 0;
      _tmp_937 <= 0;
      _tmp_938 <= 0;
      _tmp_939 <= 0;
      _tmp_940 <= 0;
      _tmp_941 <= 0;
      _tmp_942 <= 0;
      _tmp_943 <= 0;
      _tmp_944 <= 0;
      _tmp_945 <= 0;
      _tmp_946 <= 0;
      _tmp_947 <= 0;
      _tmp_948 <= 0;
      _tmp_949 <= 0;
      _tmp_950 <= 0;
      _add_tree_16_busy_reg <= 0;
    end else begin
      if(_add_tree_16_stream_oready) begin
        _add_tree_16_var0_source_ram_renable <= 0;
        _add_tree_16_var0_source_fifo_deq <= 0;
      end 
      _add_tree_16_var0_idle <= _add_tree_16_var0_idle;
      if(_add_tree_16_stream_oready) begin
        _add_tree_16_var1_source_ram_renable <= 0;
        _add_tree_16_var1_source_fifo_deq <= 0;
      end 
      _add_tree_16_var1_idle <= _add_tree_16_var1_idle;
      if(_add_tree_16_stream_oready) begin
        _add_tree_16_var2_source_ram_renable <= 0;
        _add_tree_16_var2_source_fifo_deq <= 0;
      end 
      _add_tree_16_var2_idle <= _add_tree_16_var2_idle;
      if(_add_tree_16_stream_oready) begin
        _add_tree_16_var3_source_ram_renable <= 0;
        _add_tree_16_var3_source_fifo_deq <= 0;
      end 
      _add_tree_16_var3_idle <= _add_tree_16_var3_idle;
      if(_add_tree_16_stream_oready) begin
        _add_tree_16_var4_source_ram_renable <= 0;
        _add_tree_16_var4_source_fifo_deq <= 0;
      end 
      _add_tree_16_var4_idle <= _add_tree_16_var4_idle;
      if(_add_tree_16_stream_oready) begin
        _add_tree_16_var5_source_ram_renable <= 0;
        _add_tree_16_var5_source_fifo_deq <= 0;
      end 
      _add_tree_16_var5_idle <= _add_tree_16_var5_idle;
      if(_add_tree_16_stream_oready) begin
        _add_tree_16_var6_source_ram_renable <= 0;
        _add_tree_16_var6_source_fifo_deq <= 0;
      end 
      _add_tree_16_var6_idle <= _add_tree_16_var6_idle;
      if(_add_tree_16_stream_oready) begin
        _add_tree_16_var7_source_ram_renable <= 0;
        _add_tree_16_var7_source_fifo_deq <= 0;
      end 
      _add_tree_16_var7_idle <= _add_tree_16_var7_idle;
      if(_add_tree_16_stream_oready) begin
        _add_tree_16_var8_source_ram_renable <= 0;
        _add_tree_16_var8_source_fifo_deq <= 0;
      end 
      _add_tree_16_var8_idle <= _add_tree_16_var8_idle;
      if(_add_tree_16_stream_oready) begin
        _add_tree_16_sum_sink_wenable <= 0;
        _add_tree_16_sum_sink_fifo_enq <= 0;
      end 
      if(_add_tree_16_stream_oready) begin
        __add_tree_16_stream_ivalid_1 <= _add_tree_16_stream_ivalid;
      end 
      if(_add_tree_16_stream_oready) begin
        __add_tree_16_stream_ivalid_2 <= __add_tree_16_stream_ivalid_1;
      end 
      if(_add_tree_16_stream_oready) begin
        __plusn_data_1314 <= add_tree_16_var0_data + add_tree_16_var1_data + add_tree_16_var2_data;
      end 
      if(_add_tree_16_stream_oready) begin
        __plusn_data_1315 <= add_tree_16_var3_data + add_tree_16_var4_data + add_tree_16_var5_data;
      end 
      if(_add_tree_16_stream_oready) begin
        __plusn_data_1316 <= add_tree_16_var6_data + add_tree_16_var7_data + add_tree_16_var8_data;
      end 
      if(_add_tree_16_stream_oready) begin
        __plusn_data_1317 <= __plusn_data_1314 + __plusn_data_1315 + __plusn_data_1316;
      end 
      if(__stream_conv2d_4_stream_ivalid_10 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_1304 <= __substreamoutput_data_1944;
      end 
      if(__stream_conv2d_4_stream_ivalid_10 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_1305 <= __substreamoutput_data_1963;
      end 
      if(__stream_conv2d_4_stream_ivalid_10 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_1306 <= __substreamoutput_data_1982;
      end 
      if(__stream_conv2d_4_stream_ivalid_10 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_1307 <= __substreamoutput_data_2001;
      end 
      if(__stream_conv2d_4_stream_ivalid_10 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_1308 <= __substreamoutput_data_2020;
      end 
      if(__stream_conv2d_4_stream_ivalid_10 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_1309 <= __substreamoutput_data_2039;
      end 
      if(__stream_conv2d_4_stream_ivalid_10 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_1310 <= __substreamoutput_data_2058;
      end 
      if(__stream_conv2d_4_stream_ivalid_10 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_1311 <= __substreamoutput_data_2077;
      end 
      if(__stream_conv2d_4_stream_ivalid_10 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_1312 <= __substreamoutput_data_2096;
      end 
      if(_add_tree_16_stream_oready) begin
        _tmp_935 <= _add_tree_16_source_start;
      end 
      if(_add_tree_16_stream_oready) begin
        _tmp_936 <= _tmp_935;
      end 
      if(_add_tree_16_stream_oready) begin
        _tmp_937 <= _tmp_936;
      end 
      if(_add_tree_16_stream_oready) begin
        _tmp_938 <= _add_tree_16_source_start;
      end 
      if(_add_tree_16_stream_oready) begin
        _tmp_939 <= _tmp_938;
      end 
      if(_add_tree_16_stream_oready) begin
        _tmp_940 <= _tmp_939;
      end 
      if(_add_tree_16_stream_oready) begin
        _tmp_941 <= _tmp_940;
      end 
      if(_add_tree_16_stream_oready) begin
        _tmp_942 <= _add_tree_16_source_stop;
      end 
      if(_add_tree_16_stream_oready) begin
        _tmp_943 <= _tmp_942;
      end 
      if(_add_tree_16_stream_oready) begin
        _tmp_944 <= _tmp_943;
      end 
      if(_add_tree_16_stream_oready) begin
        _tmp_945 <= _tmp_944;
      end 
      if(_add_tree_16_stream_oready) begin
        _tmp_946 <= _add_tree_16_source_busy;
      end 
      if(_add_tree_16_stream_oready) begin
        _tmp_947 <= _tmp_946;
      end 
      if(_add_tree_16_stream_oready) begin
        _tmp_948 <= _tmp_947;
      end 
      if(_add_tree_16_stream_oready) begin
        _tmp_949 <= _tmp_948;
      end 
      if(_add_tree_16_stream_oready) begin
        _tmp_950 <= _add_tree_16_sink_busy;
      end 
      if(!_add_tree_16_sink_busy && _tmp_950) begin
        _add_tree_16_busy_reg <= 0;
      end 
      if(_add_tree_16_source_busy) begin
        _add_tree_16_busy_reg <= 1;
      end 
    end
  end

  localparam _add_tree_16_fsm_1 = 1;
  localparam _add_tree_16_fsm_2 = 2;
  localparam _add_tree_16_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _add_tree_16_fsm <= _add_tree_16_fsm_init;
      _add_tree_16_source_start <= 0;
      _add_tree_16_source_busy <= 0;
      _add_tree_16_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_10 && _stream_conv2d_4_stream_oready) begin
        _add_tree_16_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _add_tree_16_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_add_tree_16_stream_oready && _tmp_937) begin
        _add_tree_16_stream_ivalid <= 1;
      end 
      if(_add_tree_16_stream_oready && 1'd0) begin
        _add_tree_16_stream_ivalid <= 0;
      end 
      case(_add_tree_16_fsm)
        _add_tree_16_fsm_init: begin
          if(_add_tree_16_run_flag) begin
            _add_tree_16_source_start <= 1;
          end 
          if(_add_tree_16_run_flag) begin
            _add_tree_16_fsm <= _add_tree_16_fsm_1;
          end 
        end
        _add_tree_16_fsm_1: begin
          if(_add_tree_16_source_start && _add_tree_16_stream_oready) begin
            _add_tree_16_source_start <= 0;
            _add_tree_16_source_busy <= 1;
          end 
          if(_add_tree_16_source_start && _add_tree_16_stream_oready) begin
            _add_tree_16_fsm <= _add_tree_16_fsm_2;
          end 
        end
        _add_tree_16_fsm_2: begin
          if(_add_tree_16_stream_oready) begin
            _add_tree_16_fsm <= _add_tree_16_fsm_3;
          end 
        end
        _add_tree_16_fsm_3: begin
          if(_add_tree_16_stream_oready && 1'd0) begin
            _add_tree_16_source_busy <= 0;
          end 
          if(_add_tree_16_stream_oready && 1'd0 && _add_tree_16_run_flag) begin
            _add_tree_16_source_start <= 1;
          end 
          if(_add_tree_16_stream_oready && 1'd0) begin
            _add_tree_16_fsm <= _add_tree_16_fsm_init;
          end 
          if(_add_tree_16_stream_oready && 1'd0 && _add_tree_16_run_flag) begin
            _add_tree_16_fsm <= _add_tree_16_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_rshift_round_clip_17_x_source_ram_renable <= 0;
      _mul_rshift_round_clip_17_x_source_fifo_deq <= 0;
      _mul_rshift_round_clip_17_x_idle <= 1;
      _mul_rshift_round_clip_17_y_source_ram_renable <= 0;
      _mul_rshift_round_clip_17_y_source_fifo_deq <= 0;
      _mul_rshift_round_clip_17_y_idle <= 1;
      _mul_rshift_round_clip_17_rshift_source_ram_renable <= 0;
      _mul_rshift_round_clip_17_rshift_source_fifo_deq <= 0;
      _mul_rshift_round_clip_17_rshift_idle <= 1;
      _mul_rshift_round_clip_17_z_sink_wenable <= 0;
      _mul_rshift_round_clip_17_z_sink_fifo_enq <= 0;
      __mul_rshift_round_clip_17_stream_ivalid_1 <= 0;
      __mul_rshift_round_clip_17_stream_ivalid_2 <= 0;
      __mul_rshift_round_clip_17_stream_ivalid_3 <= 0;
      __mul_rshift_round_clip_17_stream_ivalid_4 <= 0;
      __mul_rshift_round_clip_17_stream_ivalid_5 <= 0;
      __mul_rshift_round_clip_17_stream_ivalid_6 <= 0;
      __mul_rshift_round_clip_17_stream_ivalid_7 <= 0;
      __mul_rshift_round_clip_17_stream_ivalid_8 <= 0;
      _times_mul_odata_reg_1321 <= 0;
      __delay_data_2116_sll_1327 <= 0;
      __delay_data_2120__variable_1320 <= 0;
      __delay_data_2124_eq_1339 <= 0;
      __delay_data_2117__delay_2116_sll_1327 <= 0;
      __delay_data_2121__delay_2120__variable_1320 <= 0;
      __delay_data_2125__delay_2124_eq_1339 <= 0;
      __delay_data_2118__delay_2117__delay_2116_sll_1327 <= 0;
      __delay_data_2122__delay_2121__delay_2120__variable_1320 <= 0;
      __delay_data_2126__delay_2125__delay_2124_eq_1339 <= 0;
      __delay_data_2119__delay_2118__delay_2117__delay_2116_sll_1327 <= 0;
      __delay_data_2123__delay_2122__delay_2121____variable_1320 <= 0;
      __delay_data_2127__delay_2126__delay_2125__delay_2124_eq_1339 <= 0;
      _cond_data_1340 <= 0;
      _greaterthan_data_1341 <= 0;
      _lessthan_data_1345 <= 0;
      _greatereq_data_1349 <= 0;
      __delay_data_2128_cond_1340 <= 0;
      _cond_data_1343 <= 0;
      _cond_data_1347 <= 0;
      __delay_data_2129_greatereq_1349 <= 0;
      _cond_data_1351 <= 0;
      __variable_wdata_1318 <= 0;
      __variable_wdata_1319 <= 0;
      __variable_wdata_1320 <= 0;
      _tmp_983 <= 0;
      _tmp_984 <= 0;
      _tmp_985 <= 0;
      _tmp_986 <= 0;
      _tmp_987 <= 0;
      _tmp_988 <= 0;
      _tmp_989 <= 0;
      _tmp_990 <= 0;
      _tmp_991 <= 0;
      _tmp_992 <= 0;
      _tmp_993 <= 0;
      _tmp_994 <= 0;
      _tmp_995 <= 0;
      _tmp_996 <= 0;
      _tmp_997 <= 0;
      _tmp_998 <= 0;
      _tmp_999 <= 0;
      _tmp_1000 <= 0;
      _tmp_1001 <= 0;
      _tmp_1002 <= 0;
      _tmp_1003 <= 0;
      _tmp_1004 <= 0;
      _tmp_1005 <= 0;
      _tmp_1006 <= 0;
      _tmp_1007 <= 0;
      _tmp_1008 <= 0;
      _tmp_1009 <= 0;
      _tmp_1010 <= 0;
      _tmp_1011 <= 0;
      _tmp_1012 <= 0;
      _tmp_1013 <= 0;
      _tmp_1014 <= 0;
      _tmp_1015 <= 0;
      _tmp_1016 <= 0;
      _mul_rshift_round_clip_17_busy_reg <= 0;
    end else begin
      if(_mul_rshift_round_clip_17_stream_oready) begin
        _mul_rshift_round_clip_17_x_source_ram_renable <= 0;
        _mul_rshift_round_clip_17_x_source_fifo_deq <= 0;
      end 
      _mul_rshift_round_clip_17_x_idle <= _mul_rshift_round_clip_17_x_idle;
      if(_mul_rshift_round_clip_17_stream_oready) begin
        _mul_rshift_round_clip_17_y_source_ram_renable <= 0;
        _mul_rshift_round_clip_17_y_source_fifo_deq <= 0;
      end 
      _mul_rshift_round_clip_17_y_idle <= _mul_rshift_round_clip_17_y_idle;
      if(_mul_rshift_round_clip_17_stream_oready) begin
        _mul_rshift_round_clip_17_rshift_source_ram_renable <= 0;
        _mul_rshift_round_clip_17_rshift_source_fifo_deq <= 0;
      end 
      _mul_rshift_round_clip_17_rshift_idle <= _mul_rshift_round_clip_17_rshift_idle;
      if(_mul_rshift_round_clip_17_stream_oready) begin
        _mul_rshift_round_clip_17_z_sink_wenable <= 0;
        _mul_rshift_round_clip_17_z_sink_fifo_enq <= 0;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        __mul_rshift_round_clip_17_stream_ivalid_1 <= _mul_rshift_round_clip_17_stream_ivalid;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        __mul_rshift_round_clip_17_stream_ivalid_2 <= __mul_rshift_round_clip_17_stream_ivalid_1;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        __mul_rshift_round_clip_17_stream_ivalid_3 <= __mul_rshift_round_clip_17_stream_ivalid_2;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        __mul_rshift_round_clip_17_stream_ivalid_4 <= __mul_rshift_round_clip_17_stream_ivalid_3;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        __mul_rshift_round_clip_17_stream_ivalid_5 <= __mul_rshift_round_clip_17_stream_ivalid_4;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        __mul_rshift_round_clip_17_stream_ivalid_6 <= __mul_rshift_round_clip_17_stream_ivalid_5;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        __mul_rshift_round_clip_17_stream_ivalid_7 <= __mul_rshift_round_clip_17_stream_ivalid_6;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        __mul_rshift_round_clip_17_stream_ivalid_8 <= __mul_rshift_round_clip_17_stream_ivalid_7;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        _times_mul_odata_reg_1321 <= _times_mul_odata_1321;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        __delay_data_2116_sll_1327 <= _sll_data_1327;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        __delay_data_2120__variable_1320 <= mul_rshift_round_clip_17_rshift_data;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        __delay_data_2124_eq_1339 <= _eq_data_1339;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        __delay_data_2117__delay_2116_sll_1327 <= __delay_data_2116_sll_1327;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        __delay_data_2121__delay_2120__variable_1320 <= __delay_data_2120__variable_1320;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        __delay_data_2125__delay_2124_eq_1339 <= __delay_data_2124_eq_1339;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        __delay_data_2118__delay_2117__delay_2116_sll_1327 <= __delay_data_2117__delay_2116_sll_1327;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        __delay_data_2122__delay_2121__delay_2120__variable_1320 <= __delay_data_2121__delay_2120__variable_1320;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        __delay_data_2126__delay_2125__delay_2124_eq_1339 <= __delay_data_2125__delay_2124_eq_1339;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        __delay_data_2119__delay_2118__delay_2117__delay_2116_sll_1327 <= __delay_data_2118__delay_2117__delay_2116_sll_1327;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        __delay_data_2123__delay_2122__delay_2121____variable_1320 <= __delay_data_2122__delay_2121__delay_2120__variable_1320;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        __delay_data_2127__delay_2126__delay_2125__delay_2124_eq_1339 <= __delay_data_2126__delay_2125__delay_2124_eq_1339;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        _cond_data_1340 <= (__delay_data_2127__delay_2126__delay_2125__delay_2124_eq_1339)? _times_data_1321 : _sra_data_1337;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        _greaterthan_data_1341 <= _cond_data_1340 > 16'sd32767;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        _lessthan_data_1345 <= _cond_data_1340 < -16'sd32767;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        _greatereq_data_1349 <= _cond_data_1340 >= 1'sd0;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        __delay_data_2128_cond_1340 <= _cond_data_1340;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        _cond_data_1343 <= (_greaterthan_data_1341)? 16'sd32767 : __delay_data_2128_cond_1340;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        _cond_data_1347 <= (_lessthan_data_1345)? -16'sd32767 : __delay_data_2128_cond_1340;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        __delay_data_2129_greatereq_1349 <= _greatereq_data_1349;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        _cond_data_1351 <= (__delay_data_2129_greatereq_1349)? _cond_data_1343 : _cond_data_1347;
      end 
      if(__stream_conv2d_4_stream_ivalid_20 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_1318 <= _plus_data_2114;
      end 
      if(__stream_conv2d_4_stream_ivalid_20 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_1319 <= __delay_data_2361__delay_2360__delay_2359___cond_1576;
      end 
      if(__stream_conv2d_4_stream_ivalid_20 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_1320 <= __delay_data_2380__delay_2379__delay_2378___plus_2130;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        _tmp_983 <= _mul_rshift_round_clip_17_source_start;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        _tmp_984 <= _tmp_983;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        _tmp_985 <= _tmp_984;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        _tmp_986 <= _mul_rshift_round_clip_17_source_start;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        _tmp_987 <= _tmp_986;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        _tmp_988 <= _tmp_987;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        _tmp_989 <= _tmp_988;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        _tmp_990 <= _tmp_989;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        _tmp_991 <= _tmp_990;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        _tmp_992 <= _tmp_991;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        _tmp_993 <= _tmp_992;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        _tmp_994 <= _tmp_993;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        _tmp_995 <= _tmp_994;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        _tmp_996 <= _mul_rshift_round_clip_17_source_stop;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        _tmp_997 <= _tmp_996;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        _tmp_998 <= _tmp_997;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        _tmp_999 <= _tmp_998;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        _tmp_1000 <= _tmp_999;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        _tmp_1001 <= _tmp_1000;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        _tmp_1002 <= _tmp_1001;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        _tmp_1003 <= _tmp_1002;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        _tmp_1004 <= _tmp_1003;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        _tmp_1005 <= _tmp_1004;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        _tmp_1006 <= _mul_rshift_round_clip_17_source_busy;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        _tmp_1007 <= _tmp_1006;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        _tmp_1008 <= _tmp_1007;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        _tmp_1009 <= _tmp_1008;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        _tmp_1010 <= _tmp_1009;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        _tmp_1011 <= _tmp_1010;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        _tmp_1012 <= _tmp_1011;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        _tmp_1013 <= _tmp_1012;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        _tmp_1014 <= _tmp_1013;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        _tmp_1015 <= _tmp_1014;
      end 
      if(_mul_rshift_round_clip_17_stream_oready) begin
        _tmp_1016 <= _mul_rshift_round_clip_17_sink_busy;
      end 
      if(!_mul_rshift_round_clip_17_sink_busy && _tmp_1016) begin
        _mul_rshift_round_clip_17_busy_reg <= 0;
      end 
      if(_mul_rshift_round_clip_17_source_busy) begin
        _mul_rshift_round_clip_17_busy_reg <= 1;
      end 
      if(__stream_matmul_11_stream_ivalid_18 && _stream_matmul_11_stream_oready) begin
        __variable_wdata_1318 <= _plus_data_2243;
      end 
      if(__stream_matmul_11_stream_ivalid_18 && _stream_matmul_11_stream_oready) begin
        __variable_wdata_1319 <= __delay_data_2472__delay_2471__delay_2470___cond_2184;
      end 
      if(__stream_matmul_11_stream_ivalid_18 && _stream_matmul_11_stream_oready) begin
        __variable_wdata_1320 <= __delay_data_2489__delay_2488__delay_2487___plus_2245;
      end 
    end
  end

  localparam _mul_rshift_round_clip_17_fsm_1 = 1;
  localparam _mul_rshift_round_clip_17_fsm_2 = 2;
  localparam _mul_rshift_round_clip_17_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_rshift_round_clip_17_fsm <= _mul_rshift_round_clip_17_fsm_init;
      _mul_rshift_round_clip_17_source_start <= 0;
      _mul_rshift_round_clip_17_source_busy <= 0;
      _mul_rshift_round_clip_17_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_20 && _stream_conv2d_4_stream_oready) begin
        _mul_rshift_round_clip_17_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_rshift_round_clip_17_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_rshift_round_clip_17_stream_oready && _tmp_985) begin
        _mul_rshift_round_clip_17_stream_ivalid <= 1;
      end 
      if(_mul_rshift_round_clip_17_stream_oready && 1'd0) begin
        _mul_rshift_round_clip_17_stream_ivalid <= 0;
      end 
      if(__stream_matmul_11_stream_ivalid_18 && _stream_matmul_11_stream_oready) begin
        _mul_rshift_round_clip_17_stream_ivalid <= 1'd1;
      end 
      if(_stream_matmul_11_stream_oready && _stream_matmul_11_busy) begin
        _mul_rshift_round_clip_17_source_busy <= _stream_matmul_11_source_busy;
      end 
      case(_mul_rshift_round_clip_17_fsm)
        _mul_rshift_round_clip_17_fsm_init: begin
          if(_mul_rshift_round_clip_17_run_flag) begin
            _mul_rshift_round_clip_17_source_start <= 1;
          end 
          if(_mul_rshift_round_clip_17_run_flag) begin
            _mul_rshift_round_clip_17_fsm <= _mul_rshift_round_clip_17_fsm_1;
          end 
        end
        _mul_rshift_round_clip_17_fsm_1: begin
          if(_mul_rshift_round_clip_17_source_start && _mul_rshift_round_clip_17_stream_oready) begin
            _mul_rshift_round_clip_17_source_start <= 0;
            _mul_rshift_round_clip_17_source_busy <= 1;
          end 
          if(_mul_rshift_round_clip_17_source_start && _mul_rshift_round_clip_17_stream_oready) begin
            _mul_rshift_round_clip_17_fsm <= _mul_rshift_round_clip_17_fsm_2;
          end 
        end
        _mul_rshift_round_clip_17_fsm_2: begin
          if(_mul_rshift_round_clip_17_stream_oready) begin
            _mul_rshift_round_clip_17_fsm <= _mul_rshift_round_clip_17_fsm_3;
          end 
        end
        _mul_rshift_round_clip_17_fsm_3: begin
          if(_mul_rshift_round_clip_17_stream_oready && 1'd0) begin
            _mul_rshift_round_clip_17_source_busy <= 0;
          end 
          if(_mul_rshift_round_clip_17_stream_oready && 1'd0 && _mul_rshift_round_clip_17_run_flag) begin
            _mul_rshift_round_clip_17_source_start <= 1;
          end 
          if(_mul_rshift_round_clip_17_stream_oready && 1'd0) begin
            _mul_rshift_round_clip_17_fsm <= _mul_rshift_round_clip_17_fsm_init;
          end 
          if(_mul_rshift_round_clip_17_stream_oready && 1'd0 && _mul_rshift_round_clip_17_run_flag) begin
            _mul_rshift_round_clip_17_fsm <= _mul_rshift_round_clip_17_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_18_x_source_ram_renable <= 0;
      _mul_18_x_source_fifo_deq <= 0;
      _mul_18_x_idle <= 1;
      _mul_18_y_source_ram_renable <= 0;
      _mul_18_y_source_fifo_deq <= 0;
      _mul_18_y_idle <= 1;
      _mul_18_rshift_source_ram_renable <= 0;
      _mul_18_rshift_source_fifo_deq <= 0;
      _mul_18_rshift_idle <= 1;
      _mul_18_z_sink_wenable <= 0;
      _mul_18_z_sink_fifo_enq <= 0;
      __mul_18_stream_ivalid_1 <= 0;
      __mul_18_stream_ivalid_2 <= 0;
      __mul_18_stream_ivalid_3 <= 0;
      __mul_18_stream_ivalid_4 <= 0;
      __mul_18_stream_ivalid_5 <= 0;
      __mul_18_stream_ivalid_6 <= 0;
      __mul_18_stream_ivalid_7 <= 0;
      __mul_18_stream_ivalid_8 <= 0;
      _greaterthan_data_1355 <= 0;
      _minus_data_1357 <= 0;
      _greatereq_data_1368 <= 0;
      __delay_data_1930__variable_1352 <= 0;
      __delay_data_1933__variable_1353 <= 0;
      __delay_data_1936__variable_1354 <= 0;
      _sll_data_1359 <= 0;
      __delay_data_1927_greaterthan_1355 <= 0;
      __delay_data_1928_greatereq_1368 <= 0;
      __delay_data_1931__delay_1930__variable_1352 <= 0;
      __delay_data_1934__delay_1933__variable_1353 <= 0;
      __delay_data_1937__delay_1936__variable_1354 <= 0;
      _cond_data_1365 <= 0;
      __delay_data_1929__delay_1928_greatereq_1368 <= 0;
      __delay_data_1932__delay_1931__delay_1930__variable_1352 <= 0;
      __delay_data_1935__delay_1934__delay_1933__variable_1353 <= 0;
      __delay_data_1938__delay_1937__delay_1936__variable_1354 <= 0;
      __muladd_madd_odata_reg_1371 <= 0;
      __delay_data_1939__delay_1938__delay_1937____variable_1354 <= 0;
      __delay_data_1940__delay_1939__delay_1938____variable_1354 <= 0;
      __delay_data_1941__delay_1940__delay_1939____variable_1354 <= 0;
      __delay_data_1942__delay_1941__delay_1940____variable_1354 <= 0;
      _sra_data_1372 <= 0;
      __variable_wdata_1352 <= 0;
      __variable_wdata_1353 <= 0;
      __variable_wdata_1354 <= 0;
      _tmp_629 <= 0;
      _tmp_630 <= 0;
      _tmp_631 <= 0;
      _tmp_632 <= 0;
      _tmp_633 <= 0;
      _tmp_634 <= 0;
      _tmp_635 <= 0;
      _tmp_636 <= 0;
      _tmp_637 <= 0;
      _tmp_638 <= 0;
      _tmp_639 <= 0;
      _tmp_640 <= 0;
      _tmp_641 <= 0;
      _tmp_642 <= 0;
      _tmp_643 <= 0;
      _tmp_644 <= 0;
      _tmp_645 <= 0;
      _tmp_646 <= 0;
      _tmp_647 <= 0;
      _tmp_648 <= 0;
      _tmp_649 <= 0;
      _tmp_650 <= 0;
      _tmp_651 <= 0;
      _tmp_652 <= 0;
      _tmp_653 <= 0;
      _tmp_654 <= 0;
      _tmp_655 <= 0;
      _tmp_656 <= 0;
      _tmp_657 <= 0;
      _tmp_658 <= 0;
      _tmp_659 <= 0;
      _tmp_660 <= 0;
      _tmp_661 <= 0;
      _tmp_662 <= 0;
      _mul_18_busy_reg <= 0;
    end else begin
      if(_mul_18_stream_oready) begin
        _mul_18_x_source_ram_renable <= 0;
        _mul_18_x_source_fifo_deq <= 0;
      end 
      _mul_18_x_idle <= _mul_18_x_idle;
      if(_mul_18_stream_oready) begin
        _mul_18_y_source_ram_renable <= 0;
        _mul_18_y_source_fifo_deq <= 0;
      end 
      _mul_18_y_idle <= _mul_18_y_idle;
      if(_mul_18_stream_oready) begin
        _mul_18_rshift_source_ram_renable <= 0;
        _mul_18_rshift_source_fifo_deq <= 0;
      end 
      _mul_18_rshift_idle <= _mul_18_rshift_idle;
      if(_mul_18_stream_oready) begin
        _mul_18_z_sink_wenable <= 0;
        _mul_18_z_sink_fifo_enq <= 0;
      end 
      if(_mul_18_stream_oready) begin
        __mul_18_stream_ivalid_1 <= _mul_18_stream_ivalid;
      end 
      if(_mul_18_stream_oready) begin
        __mul_18_stream_ivalid_2 <= __mul_18_stream_ivalid_1;
      end 
      if(_mul_18_stream_oready) begin
        __mul_18_stream_ivalid_3 <= __mul_18_stream_ivalid_2;
      end 
      if(_mul_18_stream_oready) begin
        __mul_18_stream_ivalid_4 <= __mul_18_stream_ivalid_3;
      end 
      if(_mul_18_stream_oready) begin
        __mul_18_stream_ivalid_5 <= __mul_18_stream_ivalid_4;
      end 
      if(_mul_18_stream_oready) begin
        __mul_18_stream_ivalid_6 <= __mul_18_stream_ivalid_5;
      end 
      if(_mul_18_stream_oready) begin
        __mul_18_stream_ivalid_7 <= __mul_18_stream_ivalid_6;
      end 
      if(_mul_18_stream_oready) begin
        __mul_18_stream_ivalid_8 <= __mul_18_stream_ivalid_7;
      end 
      if(_mul_18_stream_oready) begin
        _greaterthan_data_1355 <= mul_18_rshift_data > 1'sd0;
      end 
      if(_mul_18_stream_oready) begin
        _minus_data_1357 <= mul_18_rshift_data - 2'sd1;
      end 
      if(_mul_18_stream_oready) begin
        _greatereq_data_1368 <= mul_18_x_data >= 1'sd0;
      end 
      if(_mul_18_stream_oready) begin
        __delay_data_1930__variable_1352 <= mul_18_x_data;
      end 
      if(_mul_18_stream_oready) begin
        __delay_data_1933__variable_1353 <= mul_18_y_data;
      end 
      if(_mul_18_stream_oready) begin
        __delay_data_1936__variable_1354 <= mul_18_rshift_data;
      end 
      if(_mul_18_stream_oready) begin
        _sll_data_1359 <= 2'sd1 << _minus_data_1357;
      end 
      if(_mul_18_stream_oready) begin
        __delay_data_1927_greaterthan_1355 <= _greaterthan_data_1355;
      end 
      if(_mul_18_stream_oready) begin
        __delay_data_1928_greatereq_1368 <= _greatereq_data_1368;
      end 
      if(_mul_18_stream_oready) begin
        __delay_data_1931__delay_1930__variable_1352 <= __delay_data_1930__variable_1352;
      end 
      if(_mul_18_stream_oready) begin
        __delay_data_1934__delay_1933__variable_1353 <= __delay_data_1933__variable_1353;
      end 
      if(_mul_18_stream_oready) begin
        __delay_data_1937__delay_1936__variable_1354 <= __delay_data_1936__variable_1354;
      end 
      if(_mul_18_stream_oready) begin
        _cond_data_1365 <= (__delay_data_1927_greaterthan_1355)? _sll_data_1359 : 1'sd0;
      end 
      if(_mul_18_stream_oready) begin
        __delay_data_1929__delay_1928_greatereq_1368 <= __delay_data_1928_greatereq_1368;
      end 
      if(_mul_18_stream_oready) begin
        __delay_data_1932__delay_1931__delay_1930__variable_1352 <= __delay_data_1931__delay_1930__variable_1352;
      end 
      if(_mul_18_stream_oready) begin
        __delay_data_1935__delay_1934__delay_1933__variable_1353 <= __delay_data_1934__delay_1933__variable_1353;
      end 
      if(_mul_18_stream_oready) begin
        __delay_data_1938__delay_1937__delay_1936__variable_1354 <= __delay_data_1937__delay_1936__variable_1354;
      end 
      if(_mul_18_stream_oready) begin
        __muladd_madd_odata_reg_1371 <= __muladd_madd_odata_1371;
      end 
      if(_mul_18_stream_oready) begin
        __delay_data_1939__delay_1938__delay_1937____variable_1354 <= __delay_data_1938__delay_1937__delay_1936__variable_1354;
      end 
      if(_mul_18_stream_oready) begin
        __delay_data_1940__delay_1939__delay_1938____variable_1354 <= __delay_data_1939__delay_1938__delay_1937____variable_1354;
      end 
      if(_mul_18_stream_oready) begin
        __delay_data_1941__delay_1940__delay_1939____variable_1354 <= __delay_data_1940__delay_1939__delay_1938____variable_1354;
      end 
      if(_mul_18_stream_oready) begin
        __delay_data_1942__delay_1941__delay_1940____variable_1354 <= __delay_data_1941__delay_1940__delay_1939____variable_1354;
      end 
      if(_mul_18_stream_oready) begin
        _sra_data_1372 <= __muladd_data_1371 >>> __delay_data_1942__delay_1941__delay_1940____variable_1354;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_1352 <= _cond_data_1909;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_1353 <= __delay_data_2268_reinterpretcast_1881;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_1354 <= _plus_data_1943;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_629 <= _mul_18_source_start;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_630 <= _tmp_629;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_631 <= _tmp_630;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_632 <= _mul_18_source_start;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_633 <= _tmp_632;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_634 <= _tmp_633;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_635 <= _tmp_634;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_636 <= _tmp_635;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_637 <= _tmp_636;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_638 <= _tmp_637;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_639 <= _tmp_638;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_640 <= _tmp_639;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_641 <= _tmp_640;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_642 <= _mul_18_source_stop;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_643 <= _tmp_642;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_644 <= _tmp_643;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_645 <= _tmp_644;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_646 <= _tmp_645;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_647 <= _tmp_646;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_648 <= _tmp_647;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_649 <= _tmp_648;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_650 <= _tmp_649;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_651 <= _tmp_650;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_652 <= _mul_18_source_busy;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_653 <= _tmp_652;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_654 <= _tmp_653;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_655 <= _tmp_654;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_656 <= _tmp_655;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_657 <= _tmp_656;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_658 <= _tmp_657;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_659 <= _tmp_658;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_660 <= _tmp_659;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_661 <= _tmp_660;
      end 
      if(_mul_18_stream_oready) begin
        _tmp_662 <= _mul_18_sink_busy;
      end 
      if(!_mul_18_sink_busy && _tmp_662) begin
        _mul_18_busy_reg <= 0;
      end 
      if(_mul_18_source_busy) begin
        _mul_18_busy_reg <= 1;
      end 
      if(__stream_matmul_11_stream_ivalid_1 && _stream_matmul_11_stream_oready) begin
        __variable_wdata_1352 <= _cond_data_2233;
      end 
      if(__stream_matmul_11_stream_ivalid_1 && _stream_matmul_11_stream_oready) begin
        __variable_wdata_1353 <= __delay_data_2405_reinterpretcast_2229;
      end 
      if(__stream_matmul_11_stream_ivalid_1 && _stream_matmul_11_stream_oready) begin
        __variable_wdata_1354 <= _plus_data_2235;
      end 
    end
  end

  localparam _mul_18_fsm_1 = 1;
  localparam _mul_18_fsm_2 = 2;
  localparam _mul_18_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_18_fsm <= _mul_18_fsm_init;
      _mul_18_source_start <= 0;
      _mul_18_source_busy <= 0;
      _mul_18_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        _mul_18_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_18_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_18_stream_oready && _tmp_631) begin
        _mul_18_stream_ivalid <= 1;
      end 
      if(_mul_18_stream_oready && 1'd0) begin
        _mul_18_stream_ivalid <= 0;
      end 
      if(__stream_matmul_11_stream_ivalid_1 && _stream_matmul_11_stream_oready) begin
        _mul_18_stream_ivalid <= 1'd1;
      end 
      if(_stream_matmul_11_stream_oready && _stream_matmul_11_busy) begin
        _mul_18_source_busy <= _stream_matmul_11_source_busy;
      end 
      case(_mul_18_fsm)
        _mul_18_fsm_init: begin
          if(_mul_18_run_flag) begin
            _mul_18_source_start <= 1;
          end 
          if(_mul_18_run_flag) begin
            _mul_18_fsm <= _mul_18_fsm_1;
          end 
        end
        _mul_18_fsm_1: begin
          if(_mul_18_source_start && _mul_18_stream_oready) begin
            _mul_18_source_start <= 0;
            _mul_18_source_busy <= 1;
          end 
          if(_mul_18_source_start && _mul_18_stream_oready) begin
            _mul_18_fsm <= _mul_18_fsm_2;
          end 
        end
        _mul_18_fsm_2: begin
          if(_mul_18_stream_oready) begin
            _mul_18_fsm <= _mul_18_fsm_3;
          end 
        end
        _mul_18_fsm_3: begin
          if(_mul_18_stream_oready && 1'd0) begin
            _mul_18_source_busy <= 0;
          end 
          if(_mul_18_stream_oready && 1'd0 && _mul_18_run_flag) begin
            _mul_18_source_start <= 1;
          end 
          if(_mul_18_stream_oready && 1'd0) begin
            _mul_18_fsm <= _mul_18_fsm_init;
          end 
          if(_mul_18_stream_oready && 1'd0 && _mul_18_run_flag) begin
            _mul_18_fsm <= _mul_18_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_19_x_source_ram_renable <= 0;
      _mul_19_x_source_fifo_deq <= 0;
      _mul_19_x_idle <= 1;
      _mul_19_y_source_ram_renable <= 0;
      _mul_19_y_source_fifo_deq <= 0;
      _mul_19_y_idle <= 1;
      _mul_19_rshift_source_ram_renable <= 0;
      _mul_19_rshift_source_fifo_deq <= 0;
      _mul_19_rshift_idle <= 1;
      _mul_19_z_sink_wenable <= 0;
      _mul_19_z_sink_fifo_enq <= 0;
      __mul_19_stream_ivalid_1 <= 0;
      __mul_19_stream_ivalid_2 <= 0;
      __mul_19_stream_ivalid_3 <= 0;
      __mul_19_stream_ivalid_4 <= 0;
      __mul_19_stream_ivalid_5 <= 0;
      __mul_19_stream_ivalid_6 <= 0;
      __mul_19_stream_ivalid_7 <= 0;
      __mul_19_stream_ivalid_8 <= 0;
      _greaterthan_data_1376 <= 0;
      _minus_data_1378 <= 0;
      _greatereq_data_1389 <= 0;
      __delay_data_1949__variable_1373 <= 0;
      __delay_data_1952__variable_1374 <= 0;
      __delay_data_1955__variable_1375 <= 0;
      _sll_data_1380 <= 0;
      __delay_data_1946_greaterthan_1376 <= 0;
      __delay_data_1947_greatereq_1389 <= 0;
      __delay_data_1950__delay_1949__variable_1373 <= 0;
      __delay_data_1953__delay_1952__variable_1374 <= 0;
      __delay_data_1956__delay_1955__variable_1375 <= 0;
      _cond_data_1386 <= 0;
      __delay_data_1948__delay_1947_greatereq_1389 <= 0;
      __delay_data_1951__delay_1950__delay_1949__variable_1373 <= 0;
      __delay_data_1954__delay_1953__delay_1952__variable_1374 <= 0;
      __delay_data_1957__delay_1956__delay_1955__variable_1375 <= 0;
      __muladd_madd_odata_reg_1392 <= 0;
      __delay_data_1958__delay_1957__delay_1956____variable_1375 <= 0;
      __delay_data_1959__delay_1958__delay_1957____variable_1375 <= 0;
      __delay_data_1960__delay_1959__delay_1958____variable_1375 <= 0;
      __delay_data_1961__delay_1960__delay_1959____variable_1375 <= 0;
      _sra_data_1393 <= 0;
      __variable_wdata_1373 <= 0;
      __variable_wdata_1374 <= 0;
      __variable_wdata_1375 <= 0;
      _tmp_663 <= 0;
      _tmp_664 <= 0;
      _tmp_665 <= 0;
      _tmp_666 <= 0;
      _tmp_667 <= 0;
      _tmp_668 <= 0;
      _tmp_669 <= 0;
      _tmp_670 <= 0;
      _tmp_671 <= 0;
      _tmp_672 <= 0;
      _tmp_673 <= 0;
      _tmp_674 <= 0;
      _tmp_675 <= 0;
      _tmp_676 <= 0;
      _tmp_677 <= 0;
      _tmp_678 <= 0;
      _tmp_679 <= 0;
      _tmp_680 <= 0;
      _tmp_681 <= 0;
      _tmp_682 <= 0;
      _tmp_683 <= 0;
      _tmp_684 <= 0;
      _tmp_685 <= 0;
      _tmp_686 <= 0;
      _tmp_687 <= 0;
      _tmp_688 <= 0;
      _tmp_689 <= 0;
      _tmp_690 <= 0;
      _tmp_691 <= 0;
      _tmp_692 <= 0;
      _tmp_693 <= 0;
      _tmp_694 <= 0;
      _tmp_695 <= 0;
      _tmp_696 <= 0;
      _mul_19_busy_reg <= 0;
    end else begin
      if(_mul_19_stream_oready) begin
        _mul_19_x_source_ram_renable <= 0;
        _mul_19_x_source_fifo_deq <= 0;
      end 
      _mul_19_x_idle <= _mul_19_x_idle;
      if(_mul_19_stream_oready) begin
        _mul_19_y_source_ram_renable <= 0;
        _mul_19_y_source_fifo_deq <= 0;
      end 
      _mul_19_y_idle <= _mul_19_y_idle;
      if(_mul_19_stream_oready) begin
        _mul_19_rshift_source_ram_renable <= 0;
        _mul_19_rshift_source_fifo_deq <= 0;
      end 
      _mul_19_rshift_idle <= _mul_19_rshift_idle;
      if(_mul_19_stream_oready) begin
        _mul_19_z_sink_wenable <= 0;
        _mul_19_z_sink_fifo_enq <= 0;
      end 
      if(_mul_19_stream_oready) begin
        __mul_19_stream_ivalid_1 <= _mul_19_stream_ivalid;
      end 
      if(_mul_19_stream_oready) begin
        __mul_19_stream_ivalid_2 <= __mul_19_stream_ivalid_1;
      end 
      if(_mul_19_stream_oready) begin
        __mul_19_stream_ivalid_3 <= __mul_19_stream_ivalid_2;
      end 
      if(_mul_19_stream_oready) begin
        __mul_19_stream_ivalid_4 <= __mul_19_stream_ivalid_3;
      end 
      if(_mul_19_stream_oready) begin
        __mul_19_stream_ivalid_5 <= __mul_19_stream_ivalid_4;
      end 
      if(_mul_19_stream_oready) begin
        __mul_19_stream_ivalid_6 <= __mul_19_stream_ivalid_5;
      end 
      if(_mul_19_stream_oready) begin
        __mul_19_stream_ivalid_7 <= __mul_19_stream_ivalid_6;
      end 
      if(_mul_19_stream_oready) begin
        __mul_19_stream_ivalid_8 <= __mul_19_stream_ivalid_7;
      end 
      if(_mul_19_stream_oready) begin
        _greaterthan_data_1376 <= mul_19_rshift_data > 1'sd0;
      end 
      if(_mul_19_stream_oready) begin
        _minus_data_1378 <= mul_19_rshift_data - 2'sd1;
      end 
      if(_mul_19_stream_oready) begin
        _greatereq_data_1389 <= mul_19_x_data >= 1'sd0;
      end 
      if(_mul_19_stream_oready) begin
        __delay_data_1949__variable_1373 <= mul_19_x_data;
      end 
      if(_mul_19_stream_oready) begin
        __delay_data_1952__variable_1374 <= mul_19_y_data;
      end 
      if(_mul_19_stream_oready) begin
        __delay_data_1955__variable_1375 <= mul_19_rshift_data;
      end 
      if(_mul_19_stream_oready) begin
        _sll_data_1380 <= 2'sd1 << _minus_data_1378;
      end 
      if(_mul_19_stream_oready) begin
        __delay_data_1946_greaterthan_1376 <= _greaterthan_data_1376;
      end 
      if(_mul_19_stream_oready) begin
        __delay_data_1947_greatereq_1389 <= _greatereq_data_1389;
      end 
      if(_mul_19_stream_oready) begin
        __delay_data_1950__delay_1949__variable_1373 <= __delay_data_1949__variable_1373;
      end 
      if(_mul_19_stream_oready) begin
        __delay_data_1953__delay_1952__variable_1374 <= __delay_data_1952__variable_1374;
      end 
      if(_mul_19_stream_oready) begin
        __delay_data_1956__delay_1955__variable_1375 <= __delay_data_1955__variable_1375;
      end 
      if(_mul_19_stream_oready) begin
        _cond_data_1386 <= (__delay_data_1946_greaterthan_1376)? _sll_data_1380 : 1'sd0;
      end 
      if(_mul_19_stream_oready) begin
        __delay_data_1948__delay_1947_greatereq_1389 <= __delay_data_1947_greatereq_1389;
      end 
      if(_mul_19_stream_oready) begin
        __delay_data_1951__delay_1950__delay_1949__variable_1373 <= __delay_data_1950__delay_1949__variable_1373;
      end 
      if(_mul_19_stream_oready) begin
        __delay_data_1954__delay_1953__delay_1952__variable_1374 <= __delay_data_1953__delay_1952__variable_1374;
      end 
      if(_mul_19_stream_oready) begin
        __delay_data_1957__delay_1956__delay_1955__variable_1375 <= __delay_data_1956__delay_1955__variable_1375;
      end 
      if(_mul_19_stream_oready) begin
        __muladd_madd_odata_reg_1392 <= __muladd_madd_odata_1392;
      end 
      if(_mul_19_stream_oready) begin
        __delay_data_1958__delay_1957__delay_1956____variable_1375 <= __delay_data_1957__delay_1956__delay_1955__variable_1375;
      end 
      if(_mul_19_stream_oready) begin
        __delay_data_1959__delay_1958__delay_1957____variable_1375 <= __delay_data_1958__delay_1957__delay_1956____variable_1375;
      end 
      if(_mul_19_stream_oready) begin
        __delay_data_1960__delay_1959__delay_1958____variable_1375 <= __delay_data_1959__delay_1958__delay_1957____variable_1375;
      end 
      if(_mul_19_stream_oready) begin
        __delay_data_1961__delay_1960__delay_1959____variable_1375 <= __delay_data_1960__delay_1959__delay_1958____variable_1375;
      end 
      if(_mul_19_stream_oready) begin
        _sra_data_1393 <= __muladd_data_1392 >>> __delay_data_1961__delay_1960__delay_1959____variable_1375;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_1373 <= _cond_data_1911;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_1374 <= __delay_data_2270_reinterpretcast_1882;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_1375 <= _plus_data_1962;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_663 <= _mul_19_source_start;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_664 <= _tmp_663;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_665 <= _tmp_664;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_666 <= _mul_19_source_start;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_667 <= _tmp_666;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_668 <= _tmp_667;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_669 <= _tmp_668;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_670 <= _tmp_669;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_671 <= _tmp_670;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_672 <= _tmp_671;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_673 <= _tmp_672;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_674 <= _tmp_673;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_675 <= _tmp_674;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_676 <= _mul_19_source_stop;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_677 <= _tmp_676;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_678 <= _tmp_677;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_679 <= _tmp_678;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_680 <= _tmp_679;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_681 <= _tmp_680;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_682 <= _tmp_681;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_683 <= _tmp_682;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_684 <= _tmp_683;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_685 <= _tmp_684;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_686 <= _mul_19_source_busy;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_687 <= _tmp_686;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_688 <= _tmp_687;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_689 <= _tmp_688;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_690 <= _tmp_689;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_691 <= _tmp_690;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_692 <= _tmp_691;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_693 <= _tmp_692;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_694 <= _tmp_693;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_695 <= _tmp_694;
      end 
      if(_mul_19_stream_oready) begin
        _tmp_696 <= _mul_19_sink_busy;
      end 
      if(!_mul_19_sink_busy && _tmp_696) begin
        _mul_19_busy_reg <= 0;
      end 
      if(_mul_19_source_busy) begin
        _mul_19_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_19_fsm_1 = 1;
  localparam _mul_19_fsm_2 = 2;
  localparam _mul_19_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_19_fsm <= _mul_19_fsm_init;
      _mul_19_source_start <= 0;
      _mul_19_source_busy <= 0;
      _mul_19_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        _mul_19_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_19_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_19_stream_oready && _tmp_665) begin
        _mul_19_stream_ivalid <= 1;
      end 
      if(_mul_19_stream_oready && 1'd0) begin
        _mul_19_stream_ivalid <= 0;
      end 
      case(_mul_19_fsm)
        _mul_19_fsm_init: begin
          if(_mul_19_run_flag) begin
            _mul_19_source_start <= 1;
          end 
          if(_mul_19_run_flag) begin
            _mul_19_fsm <= _mul_19_fsm_1;
          end 
        end
        _mul_19_fsm_1: begin
          if(_mul_19_source_start && _mul_19_stream_oready) begin
            _mul_19_source_start <= 0;
            _mul_19_source_busy <= 1;
          end 
          if(_mul_19_source_start && _mul_19_stream_oready) begin
            _mul_19_fsm <= _mul_19_fsm_2;
          end 
        end
        _mul_19_fsm_2: begin
          if(_mul_19_stream_oready) begin
            _mul_19_fsm <= _mul_19_fsm_3;
          end 
        end
        _mul_19_fsm_3: begin
          if(_mul_19_stream_oready && 1'd0) begin
            _mul_19_source_busy <= 0;
          end 
          if(_mul_19_stream_oready && 1'd0 && _mul_19_run_flag) begin
            _mul_19_source_start <= 1;
          end 
          if(_mul_19_stream_oready && 1'd0) begin
            _mul_19_fsm <= _mul_19_fsm_init;
          end 
          if(_mul_19_stream_oready && 1'd0 && _mul_19_run_flag) begin
            _mul_19_fsm <= _mul_19_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_20_x_source_ram_renable <= 0;
      _mul_20_x_source_fifo_deq <= 0;
      _mul_20_x_idle <= 1;
      _mul_20_y_source_ram_renable <= 0;
      _mul_20_y_source_fifo_deq <= 0;
      _mul_20_y_idle <= 1;
      _mul_20_rshift_source_ram_renable <= 0;
      _mul_20_rshift_source_fifo_deq <= 0;
      _mul_20_rshift_idle <= 1;
      _mul_20_z_sink_wenable <= 0;
      _mul_20_z_sink_fifo_enq <= 0;
      __mul_20_stream_ivalid_1 <= 0;
      __mul_20_stream_ivalid_2 <= 0;
      __mul_20_stream_ivalid_3 <= 0;
      __mul_20_stream_ivalid_4 <= 0;
      __mul_20_stream_ivalid_5 <= 0;
      __mul_20_stream_ivalid_6 <= 0;
      __mul_20_stream_ivalid_7 <= 0;
      __mul_20_stream_ivalid_8 <= 0;
      _greaterthan_data_1397 <= 0;
      _minus_data_1399 <= 0;
      _greatereq_data_1410 <= 0;
      __delay_data_1968__variable_1394 <= 0;
      __delay_data_1971__variable_1395 <= 0;
      __delay_data_1974__variable_1396 <= 0;
      _sll_data_1401 <= 0;
      __delay_data_1965_greaterthan_1397 <= 0;
      __delay_data_1966_greatereq_1410 <= 0;
      __delay_data_1969__delay_1968__variable_1394 <= 0;
      __delay_data_1972__delay_1971__variable_1395 <= 0;
      __delay_data_1975__delay_1974__variable_1396 <= 0;
      _cond_data_1407 <= 0;
      __delay_data_1967__delay_1966_greatereq_1410 <= 0;
      __delay_data_1970__delay_1969__delay_1968__variable_1394 <= 0;
      __delay_data_1973__delay_1972__delay_1971__variable_1395 <= 0;
      __delay_data_1976__delay_1975__delay_1974__variable_1396 <= 0;
      __muladd_madd_odata_reg_1413 <= 0;
      __delay_data_1977__delay_1976__delay_1975____variable_1396 <= 0;
      __delay_data_1978__delay_1977__delay_1976____variable_1396 <= 0;
      __delay_data_1979__delay_1978__delay_1977____variable_1396 <= 0;
      __delay_data_1980__delay_1979__delay_1978____variable_1396 <= 0;
      _sra_data_1414 <= 0;
      __variable_wdata_1394 <= 0;
      __variable_wdata_1395 <= 0;
      __variable_wdata_1396 <= 0;
      _tmp_697 <= 0;
      _tmp_698 <= 0;
      _tmp_699 <= 0;
      _tmp_700 <= 0;
      _tmp_701 <= 0;
      _tmp_702 <= 0;
      _tmp_703 <= 0;
      _tmp_704 <= 0;
      _tmp_705 <= 0;
      _tmp_706 <= 0;
      _tmp_707 <= 0;
      _tmp_708 <= 0;
      _tmp_709 <= 0;
      _tmp_710 <= 0;
      _tmp_711 <= 0;
      _tmp_712 <= 0;
      _tmp_713 <= 0;
      _tmp_714 <= 0;
      _tmp_715 <= 0;
      _tmp_716 <= 0;
      _tmp_717 <= 0;
      _tmp_718 <= 0;
      _tmp_719 <= 0;
      _tmp_720 <= 0;
      _tmp_721 <= 0;
      _tmp_722 <= 0;
      _tmp_723 <= 0;
      _tmp_724 <= 0;
      _tmp_725 <= 0;
      _tmp_726 <= 0;
      _tmp_727 <= 0;
      _tmp_728 <= 0;
      _tmp_729 <= 0;
      _tmp_730 <= 0;
      _mul_20_busy_reg <= 0;
    end else begin
      if(_mul_20_stream_oready) begin
        _mul_20_x_source_ram_renable <= 0;
        _mul_20_x_source_fifo_deq <= 0;
      end 
      _mul_20_x_idle <= _mul_20_x_idle;
      if(_mul_20_stream_oready) begin
        _mul_20_y_source_ram_renable <= 0;
        _mul_20_y_source_fifo_deq <= 0;
      end 
      _mul_20_y_idle <= _mul_20_y_idle;
      if(_mul_20_stream_oready) begin
        _mul_20_rshift_source_ram_renable <= 0;
        _mul_20_rshift_source_fifo_deq <= 0;
      end 
      _mul_20_rshift_idle <= _mul_20_rshift_idle;
      if(_mul_20_stream_oready) begin
        _mul_20_z_sink_wenable <= 0;
        _mul_20_z_sink_fifo_enq <= 0;
      end 
      if(_mul_20_stream_oready) begin
        __mul_20_stream_ivalid_1 <= _mul_20_stream_ivalid;
      end 
      if(_mul_20_stream_oready) begin
        __mul_20_stream_ivalid_2 <= __mul_20_stream_ivalid_1;
      end 
      if(_mul_20_stream_oready) begin
        __mul_20_stream_ivalid_3 <= __mul_20_stream_ivalid_2;
      end 
      if(_mul_20_stream_oready) begin
        __mul_20_stream_ivalid_4 <= __mul_20_stream_ivalid_3;
      end 
      if(_mul_20_stream_oready) begin
        __mul_20_stream_ivalid_5 <= __mul_20_stream_ivalid_4;
      end 
      if(_mul_20_stream_oready) begin
        __mul_20_stream_ivalid_6 <= __mul_20_stream_ivalid_5;
      end 
      if(_mul_20_stream_oready) begin
        __mul_20_stream_ivalid_7 <= __mul_20_stream_ivalid_6;
      end 
      if(_mul_20_stream_oready) begin
        __mul_20_stream_ivalid_8 <= __mul_20_stream_ivalid_7;
      end 
      if(_mul_20_stream_oready) begin
        _greaterthan_data_1397 <= mul_20_rshift_data > 1'sd0;
      end 
      if(_mul_20_stream_oready) begin
        _minus_data_1399 <= mul_20_rshift_data - 2'sd1;
      end 
      if(_mul_20_stream_oready) begin
        _greatereq_data_1410 <= mul_20_x_data >= 1'sd0;
      end 
      if(_mul_20_stream_oready) begin
        __delay_data_1968__variable_1394 <= mul_20_x_data;
      end 
      if(_mul_20_stream_oready) begin
        __delay_data_1971__variable_1395 <= mul_20_y_data;
      end 
      if(_mul_20_stream_oready) begin
        __delay_data_1974__variable_1396 <= mul_20_rshift_data;
      end 
      if(_mul_20_stream_oready) begin
        _sll_data_1401 <= 2'sd1 << _minus_data_1399;
      end 
      if(_mul_20_stream_oready) begin
        __delay_data_1965_greaterthan_1397 <= _greaterthan_data_1397;
      end 
      if(_mul_20_stream_oready) begin
        __delay_data_1966_greatereq_1410 <= _greatereq_data_1410;
      end 
      if(_mul_20_stream_oready) begin
        __delay_data_1969__delay_1968__variable_1394 <= __delay_data_1968__variable_1394;
      end 
      if(_mul_20_stream_oready) begin
        __delay_data_1972__delay_1971__variable_1395 <= __delay_data_1971__variable_1395;
      end 
      if(_mul_20_stream_oready) begin
        __delay_data_1975__delay_1974__variable_1396 <= __delay_data_1974__variable_1396;
      end 
      if(_mul_20_stream_oready) begin
        _cond_data_1407 <= (__delay_data_1965_greaterthan_1397)? _sll_data_1401 : 1'sd0;
      end 
      if(_mul_20_stream_oready) begin
        __delay_data_1967__delay_1966_greatereq_1410 <= __delay_data_1966_greatereq_1410;
      end 
      if(_mul_20_stream_oready) begin
        __delay_data_1970__delay_1969__delay_1968__variable_1394 <= __delay_data_1969__delay_1968__variable_1394;
      end 
      if(_mul_20_stream_oready) begin
        __delay_data_1973__delay_1972__delay_1971__variable_1395 <= __delay_data_1972__delay_1971__variable_1395;
      end 
      if(_mul_20_stream_oready) begin
        __delay_data_1976__delay_1975__delay_1974__variable_1396 <= __delay_data_1975__delay_1974__variable_1396;
      end 
      if(_mul_20_stream_oready) begin
        __muladd_madd_odata_reg_1413 <= __muladd_madd_odata_1413;
      end 
      if(_mul_20_stream_oready) begin
        __delay_data_1977__delay_1976__delay_1975____variable_1396 <= __delay_data_1976__delay_1975__delay_1974__variable_1396;
      end 
      if(_mul_20_stream_oready) begin
        __delay_data_1978__delay_1977__delay_1976____variable_1396 <= __delay_data_1977__delay_1976__delay_1975____variable_1396;
      end 
      if(_mul_20_stream_oready) begin
        __delay_data_1979__delay_1978__delay_1977____variable_1396 <= __delay_data_1978__delay_1977__delay_1976____variable_1396;
      end 
      if(_mul_20_stream_oready) begin
        __delay_data_1980__delay_1979__delay_1978____variable_1396 <= __delay_data_1979__delay_1978__delay_1977____variable_1396;
      end 
      if(_mul_20_stream_oready) begin
        _sra_data_1414 <= __muladd_data_1413 >>> __delay_data_1980__delay_1979__delay_1978____variable_1396;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_1394 <= _cond_data_1913;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_1395 <= __delay_data_2272_reinterpretcast_1883;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_1396 <= _plus_data_1981;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_697 <= _mul_20_source_start;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_698 <= _tmp_697;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_699 <= _tmp_698;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_700 <= _mul_20_source_start;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_701 <= _tmp_700;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_702 <= _tmp_701;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_703 <= _tmp_702;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_704 <= _tmp_703;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_705 <= _tmp_704;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_706 <= _tmp_705;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_707 <= _tmp_706;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_708 <= _tmp_707;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_709 <= _tmp_708;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_710 <= _mul_20_source_stop;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_711 <= _tmp_710;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_712 <= _tmp_711;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_713 <= _tmp_712;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_714 <= _tmp_713;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_715 <= _tmp_714;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_716 <= _tmp_715;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_717 <= _tmp_716;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_718 <= _tmp_717;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_719 <= _tmp_718;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_720 <= _mul_20_source_busy;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_721 <= _tmp_720;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_722 <= _tmp_721;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_723 <= _tmp_722;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_724 <= _tmp_723;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_725 <= _tmp_724;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_726 <= _tmp_725;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_727 <= _tmp_726;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_728 <= _tmp_727;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_729 <= _tmp_728;
      end 
      if(_mul_20_stream_oready) begin
        _tmp_730 <= _mul_20_sink_busy;
      end 
      if(!_mul_20_sink_busy && _tmp_730) begin
        _mul_20_busy_reg <= 0;
      end 
      if(_mul_20_source_busy) begin
        _mul_20_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_20_fsm_1 = 1;
  localparam _mul_20_fsm_2 = 2;
  localparam _mul_20_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_20_fsm <= _mul_20_fsm_init;
      _mul_20_source_start <= 0;
      _mul_20_source_busy <= 0;
      _mul_20_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        _mul_20_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_20_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_20_stream_oready && _tmp_699) begin
        _mul_20_stream_ivalid <= 1;
      end 
      if(_mul_20_stream_oready && 1'd0) begin
        _mul_20_stream_ivalid <= 0;
      end 
      case(_mul_20_fsm)
        _mul_20_fsm_init: begin
          if(_mul_20_run_flag) begin
            _mul_20_source_start <= 1;
          end 
          if(_mul_20_run_flag) begin
            _mul_20_fsm <= _mul_20_fsm_1;
          end 
        end
        _mul_20_fsm_1: begin
          if(_mul_20_source_start && _mul_20_stream_oready) begin
            _mul_20_source_start <= 0;
            _mul_20_source_busy <= 1;
          end 
          if(_mul_20_source_start && _mul_20_stream_oready) begin
            _mul_20_fsm <= _mul_20_fsm_2;
          end 
        end
        _mul_20_fsm_2: begin
          if(_mul_20_stream_oready) begin
            _mul_20_fsm <= _mul_20_fsm_3;
          end 
        end
        _mul_20_fsm_3: begin
          if(_mul_20_stream_oready && 1'd0) begin
            _mul_20_source_busy <= 0;
          end 
          if(_mul_20_stream_oready && 1'd0 && _mul_20_run_flag) begin
            _mul_20_source_start <= 1;
          end 
          if(_mul_20_stream_oready && 1'd0) begin
            _mul_20_fsm <= _mul_20_fsm_init;
          end 
          if(_mul_20_stream_oready && 1'd0 && _mul_20_run_flag) begin
            _mul_20_fsm <= _mul_20_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_21_x_source_ram_renable <= 0;
      _mul_21_x_source_fifo_deq <= 0;
      _mul_21_x_idle <= 1;
      _mul_21_y_source_ram_renable <= 0;
      _mul_21_y_source_fifo_deq <= 0;
      _mul_21_y_idle <= 1;
      _mul_21_rshift_source_ram_renable <= 0;
      _mul_21_rshift_source_fifo_deq <= 0;
      _mul_21_rshift_idle <= 1;
      _mul_21_z_sink_wenable <= 0;
      _mul_21_z_sink_fifo_enq <= 0;
      __mul_21_stream_ivalid_1 <= 0;
      __mul_21_stream_ivalid_2 <= 0;
      __mul_21_stream_ivalid_3 <= 0;
      __mul_21_stream_ivalid_4 <= 0;
      __mul_21_stream_ivalid_5 <= 0;
      __mul_21_stream_ivalid_6 <= 0;
      __mul_21_stream_ivalid_7 <= 0;
      __mul_21_stream_ivalid_8 <= 0;
      _greaterthan_data_1418 <= 0;
      _minus_data_1420 <= 0;
      _greatereq_data_1431 <= 0;
      __delay_data_1987__variable_1415 <= 0;
      __delay_data_1990__variable_1416 <= 0;
      __delay_data_1993__variable_1417 <= 0;
      _sll_data_1422 <= 0;
      __delay_data_1984_greaterthan_1418 <= 0;
      __delay_data_1985_greatereq_1431 <= 0;
      __delay_data_1988__delay_1987__variable_1415 <= 0;
      __delay_data_1991__delay_1990__variable_1416 <= 0;
      __delay_data_1994__delay_1993__variable_1417 <= 0;
      _cond_data_1428 <= 0;
      __delay_data_1986__delay_1985_greatereq_1431 <= 0;
      __delay_data_1989__delay_1988__delay_1987__variable_1415 <= 0;
      __delay_data_1992__delay_1991__delay_1990__variable_1416 <= 0;
      __delay_data_1995__delay_1994__delay_1993__variable_1417 <= 0;
      __muladd_madd_odata_reg_1434 <= 0;
      __delay_data_1996__delay_1995__delay_1994____variable_1417 <= 0;
      __delay_data_1997__delay_1996__delay_1995____variable_1417 <= 0;
      __delay_data_1998__delay_1997__delay_1996____variable_1417 <= 0;
      __delay_data_1999__delay_1998__delay_1997____variable_1417 <= 0;
      _sra_data_1435 <= 0;
      __variable_wdata_1415 <= 0;
      __variable_wdata_1416 <= 0;
      __variable_wdata_1417 <= 0;
      _tmp_731 <= 0;
      _tmp_732 <= 0;
      _tmp_733 <= 0;
      _tmp_734 <= 0;
      _tmp_735 <= 0;
      _tmp_736 <= 0;
      _tmp_737 <= 0;
      _tmp_738 <= 0;
      _tmp_739 <= 0;
      _tmp_740 <= 0;
      _tmp_741 <= 0;
      _tmp_742 <= 0;
      _tmp_743 <= 0;
      _tmp_744 <= 0;
      _tmp_745 <= 0;
      _tmp_746 <= 0;
      _tmp_747 <= 0;
      _tmp_748 <= 0;
      _tmp_749 <= 0;
      _tmp_750 <= 0;
      _tmp_751 <= 0;
      _tmp_752 <= 0;
      _tmp_753 <= 0;
      _tmp_754 <= 0;
      _tmp_755 <= 0;
      _tmp_756 <= 0;
      _tmp_757 <= 0;
      _tmp_758 <= 0;
      _tmp_759 <= 0;
      _tmp_760 <= 0;
      _tmp_761 <= 0;
      _tmp_762 <= 0;
      _tmp_763 <= 0;
      _tmp_764 <= 0;
      _mul_21_busy_reg <= 0;
    end else begin
      if(_mul_21_stream_oready) begin
        _mul_21_x_source_ram_renable <= 0;
        _mul_21_x_source_fifo_deq <= 0;
      end 
      _mul_21_x_idle <= _mul_21_x_idle;
      if(_mul_21_stream_oready) begin
        _mul_21_y_source_ram_renable <= 0;
        _mul_21_y_source_fifo_deq <= 0;
      end 
      _mul_21_y_idle <= _mul_21_y_idle;
      if(_mul_21_stream_oready) begin
        _mul_21_rshift_source_ram_renable <= 0;
        _mul_21_rshift_source_fifo_deq <= 0;
      end 
      _mul_21_rshift_idle <= _mul_21_rshift_idle;
      if(_mul_21_stream_oready) begin
        _mul_21_z_sink_wenable <= 0;
        _mul_21_z_sink_fifo_enq <= 0;
      end 
      if(_mul_21_stream_oready) begin
        __mul_21_stream_ivalid_1 <= _mul_21_stream_ivalid;
      end 
      if(_mul_21_stream_oready) begin
        __mul_21_stream_ivalid_2 <= __mul_21_stream_ivalid_1;
      end 
      if(_mul_21_stream_oready) begin
        __mul_21_stream_ivalid_3 <= __mul_21_stream_ivalid_2;
      end 
      if(_mul_21_stream_oready) begin
        __mul_21_stream_ivalid_4 <= __mul_21_stream_ivalid_3;
      end 
      if(_mul_21_stream_oready) begin
        __mul_21_stream_ivalid_5 <= __mul_21_stream_ivalid_4;
      end 
      if(_mul_21_stream_oready) begin
        __mul_21_stream_ivalid_6 <= __mul_21_stream_ivalid_5;
      end 
      if(_mul_21_stream_oready) begin
        __mul_21_stream_ivalid_7 <= __mul_21_stream_ivalid_6;
      end 
      if(_mul_21_stream_oready) begin
        __mul_21_stream_ivalid_8 <= __mul_21_stream_ivalid_7;
      end 
      if(_mul_21_stream_oready) begin
        _greaterthan_data_1418 <= mul_21_rshift_data > 1'sd0;
      end 
      if(_mul_21_stream_oready) begin
        _minus_data_1420 <= mul_21_rshift_data - 2'sd1;
      end 
      if(_mul_21_stream_oready) begin
        _greatereq_data_1431 <= mul_21_x_data >= 1'sd0;
      end 
      if(_mul_21_stream_oready) begin
        __delay_data_1987__variable_1415 <= mul_21_x_data;
      end 
      if(_mul_21_stream_oready) begin
        __delay_data_1990__variable_1416 <= mul_21_y_data;
      end 
      if(_mul_21_stream_oready) begin
        __delay_data_1993__variable_1417 <= mul_21_rshift_data;
      end 
      if(_mul_21_stream_oready) begin
        _sll_data_1422 <= 2'sd1 << _minus_data_1420;
      end 
      if(_mul_21_stream_oready) begin
        __delay_data_1984_greaterthan_1418 <= _greaterthan_data_1418;
      end 
      if(_mul_21_stream_oready) begin
        __delay_data_1985_greatereq_1431 <= _greatereq_data_1431;
      end 
      if(_mul_21_stream_oready) begin
        __delay_data_1988__delay_1987__variable_1415 <= __delay_data_1987__variable_1415;
      end 
      if(_mul_21_stream_oready) begin
        __delay_data_1991__delay_1990__variable_1416 <= __delay_data_1990__variable_1416;
      end 
      if(_mul_21_stream_oready) begin
        __delay_data_1994__delay_1993__variable_1417 <= __delay_data_1993__variable_1417;
      end 
      if(_mul_21_stream_oready) begin
        _cond_data_1428 <= (__delay_data_1984_greaterthan_1418)? _sll_data_1422 : 1'sd0;
      end 
      if(_mul_21_stream_oready) begin
        __delay_data_1986__delay_1985_greatereq_1431 <= __delay_data_1985_greatereq_1431;
      end 
      if(_mul_21_stream_oready) begin
        __delay_data_1989__delay_1988__delay_1987__variable_1415 <= __delay_data_1988__delay_1987__variable_1415;
      end 
      if(_mul_21_stream_oready) begin
        __delay_data_1992__delay_1991__delay_1990__variable_1416 <= __delay_data_1991__delay_1990__variable_1416;
      end 
      if(_mul_21_stream_oready) begin
        __delay_data_1995__delay_1994__delay_1993__variable_1417 <= __delay_data_1994__delay_1993__variable_1417;
      end 
      if(_mul_21_stream_oready) begin
        __muladd_madd_odata_reg_1434 <= __muladd_madd_odata_1434;
      end 
      if(_mul_21_stream_oready) begin
        __delay_data_1996__delay_1995__delay_1994____variable_1417 <= __delay_data_1995__delay_1994__delay_1993__variable_1417;
      end 
      if(_mul_21_stream_oready) begin
        __delay_data_1997__delay_1996__delay_1995____variable_1417 <= __delay_data_1996__delay_1995__delay_1994____variable_1417;
      end 
      if(_mul_21_stream_oready) begin
        __delay_data_1998__delay_1997__delay_1996____variable_1417 <= __delay_data_1997__delay_1996__delay_1995____variable_1417;
      end 
      if(_mul_21_stream_oready) begin
        __delay_data_1999__delay_1998__delay_1997____variable_1417 <= __delay_data_1998__delay_1997__delay_1996____variable_1417;
      end 
      if(_mul_21_stream_oready) begin
        _sra_data_1435 <= __muladd_data_1434 >>> __delay_data_1999__delay_1998__delay_1997____variable_1417;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_1415 <= _cond_data_1915;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_1416 <= __delay_data_2274_reinterpretcast_1884;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_1417 <= _plus_data_2000;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_731 <= _mul_21_source_start;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_732 <= _tmp_731;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_733 <= _tmp_732;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_734 <= _mul_21_source_start;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_735 <= _tmp_734;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_736 <= _tmp_735;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_737 <= _tmp_736;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_738 <= _tmp_737;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_739 <= _tmp_738;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_740 <= _tmp_739;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_741 <= _tmp_740;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_742 <= _tmp_741;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_743 <= _tmp_742;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_744 <= _mul_21_source_stop;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_745 <= _tmp_744;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_746 <= _tmp_745;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_747 <= _tmp_746;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_748 <= _tmp_747;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_749 <= _tmp_748;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_750 <= _tmp_749;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_751 <= _tmp_750;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_752 <= _tmp_751;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_753 <= _tmp_752;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_754 <= _mul_21_source_busy;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_755 <= _tmp_754;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_756 <= _tmp_755;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_757 <= _tmp_756;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_758 <= _tmp_757;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_759 <= _tmp_758;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_760 <= _tmp_759;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_761 <= _tmp_760;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_762 <= _tmp_761;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_763 <= _tmp_762;
      end 
      if(_mul_21_stream_oready) begin
        _tmp_764 <= _mul_21_sink_busy;
      end 
      if(!_mul_21_sink_busy && _tmp_764) begin
        _mul_21_busy_reg <= 0;
      end 
      if(_mul_21_source_busy) begin
        _mul_21_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_21_fsm_1 = 1;
  localparam _mul_21_fsm_2 = 2;
  localparam _mul_21_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_21_fsm <= _mul_21_fsm_init;
      _mul_21_source_start <= 0;
      _mul_21_source_busy <= 0;
      _mul_21_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        _mul_21_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_21_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_21_stream_oready && _tmp_733) begin
        _mul_21_stream_ivalid <= 1;
      end 
      if(_mul_21_stream_oready && 1'd0) begin
        _mul_21_stream_ivalid <= 0;
      end 
      case(_mul_21_fsm)
        _mul_21_fsm_init: begin
          if(_mul_21_run_flag) begin
            _mul_21_source_start <= 1;
          end 
          if(_mul_21_run_flag) begin
            _mul_21_fsm <= _mul_21_fsm_1;
          end 
        end
        _mul_21_fsm_1: begin
          if(_mul_21_source_start && _mul_21_stream_oready) begin
            _mul_21_source_start <= 0;
            _mul_21_source_busy <= 1;
          end 
          if(_mul_21_source_start && _mul_21_stream_oready) begin
            _mul_21_fsm <= _mul_21_fsm_2;
          end 
        end
        _mul_21_fsm_2: begin
          if(_mul_21_stream_oready) begin
            _mul_21_fsm <= _mul_21_fsm_3;
          end 
        end
        _mul_21_fsm_3: begin
          if(_mul_21_stream_oready && 1'd0) begin
            _mul_21_source_busy <= 0;
          end 
          if(_mul_21_stream_oready && 1'd0 && _mul_21_run_flag) begin
            _mul_21_source_start <= 1;
          end 
          if(_mul_21_stream_oready && 1'd0) begin
            _mul_21_fsm <= _mul_21_fsm_init;
          end 
          if(_mul_21_stream_oready && 1'd0 && _mul_21_run_flag) begin
            _mul_21_fsm <= _mul_21_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_22_x_source_ram_renable <= 0;
      _mul_22_x_source_fifo_deq <= 0;
      _mul_22_x_idle <= 1;
      _mul_22_y_source_ram_renable <= 0;
      _mul_22_y_source_fifo_deq <= 0;
      _mul_22_y_idle <= 1;
      _mul_22_rshift_source_ram_renable <= 0;
      _mul_22_rshift_source_fifo_deq <= 0;
      _mul_22_rshift_idle <= 1;
      _mul_22_z_sink_wenable <= 0;
      _mul_22_z_sink_fifo_enq <= 0;
      __mul_22_stream_ivalid_1 <= 0;
      __mul_22_stream_ivalid_2 <= 0;
      __mul_22_stream_ivalid_3 <= 0;
      __mul_22_stream_ivalid_4 <= 0;
      __mul_22_stream_ivalid_5 <= 0;
      __mul_22_stream_ivalid_6 <= 0;
      __mul_22_stream_ivalid_7 <= 0;
      __mul_22_stream_ivalid_8 <= 0;
      _greaterthan_data_1439 <= 0;
      _minus_data_1441 <= 0;
      _greatereq_data_1452 <= 0;
      __delay_data_2006__variable_1436 <= 0;
      __delay_data_2009__variable_1437 <= 0;
      __delay_data_2012__variable_1438 <= 0;
      _sll_data_1443 <= 0;
      __delay_data_2003_greaterthan_1439 <= 0;
      __delay_data_2004_greatereq_1452 <= 0;
      __delay_data_2007__delay_2006__variable_1436 <= 0;
      __delay_data_2010__delay_2009__variable_1437 <= 0;
      __delay_data_2013__delay_2012__variable_1438 <= 0;
      _cond_data_1449 <= 0;
      __delay_data_2005__delay_2004_greatereq_1452 <= 0;
      __delay_data_2008__delay_2007__delay_2006__variable_1436 <= 0;
      __delay_data_2011__delay_2010__delay_2009__variable_1437 <= 0;
      __delay_data_2014__delay_2013__delay_2012__variable_1438 <= 0;
      __muladd_madd_odata_reg_1455 <= 0;
      __delay_data_2015__delay_2014__delay_2013____variable_1438 <= 0;
      __delay_data_2016__delay_2015__delay_2014____variable_1438 <= 0;
      __delay_data_2017__delay_2016__delay_2015____variable_1438 <= 0;
      __delay_data_2018__delay_2017__delay_2016____variable_1438 <= 0;
      _sra_data_1456 <= 0;
      __variable_wdata_1436 <= 0;
      __variable_wdata_1437 <= 0;
      __variable_wdata_1438 <= 0;
      _tmp_765 <= 0;
      _tmp_766 <= 0;
      _tmp_767 <= 0;
      _tmp_768 <= 0;
      _tmp_769 <= 0;
      _tmp_770 <= 0;
      _tmp_771 <= 0;
      _tmp_772 <= 0;
      _tmp_773 <= 0;
      _tmp_774 <= 0;
      _tmp_775 <= 0;
      _tmp_776 <= 0;
      _tmp_777 <= 0;
      _tmp_778 <= 0;
      _tmp_779 <= 0;
      _tmp_780 <= 0;
      _tmp_781 <= 0;
      _tmp_782 <= 0;
      _tmp_783 <= 0;
      _tmp_784 <= 0;
      _tmp_785 <= 0;
      _tmp_786 <= 0;
      _tmp_787 <= 0;
      _tmp_788 <= 0;
      _tmp_789 <= 0;
      _tmp_790 <= 0;
      _tmp_791 <= 0;
      _tmp_792 <= 0;
      _tmp_793 <= 0;
      _tmp_794 <= 0;
      _tmp_795 <= 0;
      _tmp_796 <= 0;
      _tmp_797 <= 0;
      _tmp_798 <= 0;
      _mul_22_busy_reg <= 0;
    end else begin
      if(_mul_22_stream_oready) begin
        _mul_22_x_source_ram_renable <= 0;
        _mul_22_x_source_fifo_deq <= 0;
      end 
      _mul_22_x_idle <= _mul_22_x_idle;
      if(_mul_22_stream_oready) begin
        _mul_22_y_source_ram_renable <= 0;
        _mul_22_y_source_fifo_deq <= 0;
      end 
      _mul_22_y_idle <= _mul_22_y_idle;
      if(_mul_22_stream_oready) begin
        _mul_22_rshift_source_ram_renable <= 0;
        _mul_22_rshift_source_fifo_deq <= 0;
      end 
      _mul_22_rshift_idle <= _mul_22_rshift_idle;
      if(_mul_22_stream_oready) begin
        _mul_22_z_sink_wenable <= 0;
        _mul_22_z_sink_fifo_enq <= 0;
      end 
      if(_mul_22_stream_oready) begin
        __mul_22_stream_ivalid_1 <= _mul_22_stream_ivalid;
      end 
      if(_mul_22_stream_oready) begin
        __mul_22_stream_ivalid_2 <= __mul_22_stream_ivalid_1;
      end 
      if(_mul_22_stream_oready) begin
        __mul_22_stream_ivalid_3 <= __mul_22_stream_ivalid_2;
      end 
      if(_mul_22_stream_oready) begin
        __mul_22_stream_ivalid_4 <= __mul_22_stream_ivalid_3;
      end 
      if(_mul_22_stream_oready) begin
        __mul_22_stream_ivalid_5 <= __mul_22_stream_ivalid_4;
      end 
      if(_mul_22_stream_oready) begin
        __mul_22_stream_ivalid_6 <= __mul_22_stream_ivalid_5;
      end 
      if(_mul_22_stream_oready) begin
        __mul_22_stream_ivalid_7 <= __mul_22_stream_ivalid_6;
      end 
      if(_mul_22_stream_oready) begin
        __mul_22_stream_ivalid_8 <= __mul_22_stream_ivalid_7;
      end 
      if(_mul_22_stream_oready) begin
        _greaterthan_data_1439 <= mul_22_rshift_data > 1'sd0;
      end 
      if(_mul_22_stream_oready) begin
        _minus_data_1441 <= mul_22_rshift_data - 2'sd1;
      end 
      if(_mul_22_stream_oready) begin
        _greatereq_data_1452 <= mul_22_x_data >= 1'sd0;
      end 
      if(_mul_22_stream_oready) begin
        __delay_data_2006__variable_1436 <= mul_22_x_data;
      end 
      if(_mul_22_stream_oready) begin
        __delay_data_2009__variable_1437 <= mul_22_y_data;
      end 
      if(_mul_22_stream_oready) begin
        __delay_data_2012__variable_1438 <= mul_22_rshift_data;
      end 
      if(_mul_22_stream_oready) begin
        _sll_data_1443 <= 2'sd1 << _minus_data_1441;
      end 
      if(_mul_22_stream_oready) begin
        __delay_data_2003_greaterthan_1439 <= _greaterthan_data_1439;
      end 
      if(_mul_22_stream_oready) begin
        __delay_data_2004_greatereq_1452 <= _greatereq_data_1452;
      end 
      if(_mul_22_stream_oready) begin
        __delay_data_2007__delay_2006__variable_1436 <= __delay_data_2006__variable_1436;
      end 
      if(_mul_22_stream_oready) begin
        __delay_data_2010__delay_2009__variable_1437 <= __delay_data_2009__variable_1437;
      end 
      if(_mul_22_stream_oready) begin
        __delay_data_2013__delay_2012__variable_1438 <= __delay_data_2012__variable_1438;
      end 
      if(_mul_22_stream_oready) begin
        _cond_data_1449 <= (__delay_data_2003_greaterthan_1439)? _sll_data_1443 : 1'sd0;
      end 
      if(_mul_22_stream_oready) begin
        __delay_data_2005__delay_2004_greatereq_1452 <= __delay_data_2004_greatereq_1452;
      end 
      if(_mul_22_stream_oready) begin
        __delay_data_2008__delay_2007__delay_2006__variable_1436 <= __delay_data_2007__delay_2006__variable_1436;
      end 
      if(_mul_22_stream_oready) begin
        __delay_data_2011__delay_2010__delay_2009__variable_1437 <= __delay_data_2010__delay_2009__variable_1437;
      end 
      if(_mul_22_stream_oready) begin
        __delay_data_2014__delay_2013__delay_2012__variable_1438 <= __delay_data_2013__delay_2012__variable_1438;
      end 
      if(_mul_22_stream_oready) begin
        __muladd_madd_odata_reg_1455 <= __muladd_madd_odata_1455;
      end 
      if(_mul_22_stream_oready) begin
        __delay_data_2015__delay_2014__delay_2013____variable_1438 <= __delay_data_2014__delay_2013__delay_2012__variable_1438;
      end 
      if(_mul_22_stream_oready) begin
        __delay_data_2016__delay_2015__delay_2014____variable_1438 <= __delay_data_2015__delay_2014__delay_2013____variable_1438;
      end 
      if(_mul_22_stream_oready) begin
        __delay_data_2017__delay_2016__delay_2015____variable_1438 <= __delay_data_2016__delay_2015__delay_2014____variable_1438;
      end 
      if(_mul_22_stream_oready) begin
        __delay_data_2018__delay_2017__delay_2016____variable_1438 <= __delay_data_2017__delay_2016__delay_2015____variable_1438;
      end 
      if(_mul_22_stream_oready) begin
        _sra_data_1456 <= __muladd_data_1455 >>> __delay_data_2018__delay_2017__delay_2016____variable_1438;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_1436 <= _cond_data_1917;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_1437 <= __delay_data_2276_reinterpretcast_1885;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_1438 <= _plus_data_2019;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_765 <= _mul_22_source_start;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_766 <= _tmp_765;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_767 <= _tmp_766;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_768 <= _mul_22_source_start;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_769 <= _tmp_768;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_770 <= _tmp_769;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_771 <= _tmp_770;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_772 <= _tmp_771;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_773 <= _tmp_772;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_774 <= _tmp_773;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_775 <= _tmp_774;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_776 <= _tmp_775;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_777 <= _tmp_776;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_778 <= _mul_22_source_stop;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_779 <= _tmp_778;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_780 <= _tmp_779;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_781 <= _tmp_780;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_782 <= _tmp_781;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_783 <= _tmp_782;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_784 <= _tmp_783;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_785 <= _tmp_784;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_786 <= _tmp_785;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_787 <= _tmp_786;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_788 <= _mul_22_source_busy;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_789 <= _tmp_788;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_790 <= _tmp_789;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_791 <= _tmp_790;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_792 <= _tmp_791;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_793 <= _tmp_792;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_794 <= _tmp_793;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_795 <= _tmp_794;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_796 <= _tmp_795;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_797 <= _tmp_796;
      end 
      if(_mul_22_stream_oready) begin
        _tmp_798 <= _mul_22_sink_busy;
      end 
      if(!_mul_22_sink_busy && _tmp_798) begin
        _mul_22_busy_reg <= 0;
      end 
      if(_mul_22_source_busy) begin
        _mul_22_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_22_fsm_1 = 1;
  localparam _mul_22_fsm_2 = 2;
  localparam _mul_22_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_22_fsm <= _mul_22_fsm_init;
      _mul_22_source_start <= 0;
      _mul_22_source_busy <= 0;
      _mul_22_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        _mul_22_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_22_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_22_stream_oready && _tmp_767) begin
        _mul_22_stream_ivalid <= 1;
      end 
      if(_mul_22_stream_oready && 1'd0) begin
        _mul_22_stream_ivalid <= 0;
      end 
      case(_mul_22_fsm)
        _mul_22_fsm_init: begin
          if(_mul_22_run_flag) begin
            _mul_22_source_start <= 1;
          end 
          if(_mul_22_run_flag) begin
            _mul_22_fsm <= _mul_22_fsm_1;
          end 
        end
        _mul_22_fsm_1: begin
          if(_mul_22_source_start && _mul_22_stream_oready) begin
            _mul_22_source_start <= 0;
            _mul_22_source_busy <= 1;
          end 
          if(_mul_22_source_start && _mul_22_stream_oready) begin
            _mul_22_fsm <= _mul_22_fsm_2;
          end 
        end
        _mul_22_fsm_2: begin
          if(_mul_22_stream_oready) begin
            _mul_22_fsm <= _mul_22_fsm_3;
          end 
        end
        _mul_22_fsm_3: begin
          if(_mul_22_stream_oready && 1'd0) begin
            _mul_22_source_busy <= 0;
          end 
          if(_mul_22_stream_oready && 1'd0 && _mul_22_run_flag) begin
            _mul_22_source_start <= 1;
          end 
          if(_mul_22_stream_oready && 1'd0) begin
            _mul_22_fsm <= _mul_22_fsm_init;
          end 
          if(_mul_22_stream_oready && 1'd0 && _mul_22_run_flag) begin
            _mul_22_fsm <= _mul_22_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_23_x_source_ram_renable <= 0;
      _mul_23_x_source_fifo_deq <= 0;
      _mul_23_x_idle <= 1;
      _mul_23_y_source_ram_renable <= 0;
      _mul_23_y_source_fifo_deq <= 0;
      _mul_23_y_idle <= 1;
      _mul_23_rshift_source_ram_renable <= 0;
      _mul_23_rshift_source_fifo_deq <= 0;
      _mul_23_rshift_idle <= 1;
      _mul_23_z_sink_wenable <= 0;
      _mul_23_z_sink_fifo_enq <= 0;
      __mul_23_stream_ivalid_1 <= 0;
      __mul_23_stream_ivalid_2 <= 0;
      __mul_23_stream_ivalid_3 <= 0;
      __mul_23_stream_ivalid_4 <= 0;
      __mul_23_stream_ivalid_5 <= 0;
      __mul_23_stream_ivalid_6 <= 0;
      __mul_23_stream_ivalid_7 <= 0;
      __mul_23_stream_ivalid_8 <= 0;
      _greaterthan_data_1460 <= 0;
      _minus_data_1462 <= 0;
      _greatereq_data_1473 <= 0;
      __delay_data_2025__variable_1457 <= 0;
      __delay_data_2028__variable_1458 <= 0;
      __delay_data_2031__variable_1459 <= 0;
      _sll_data_1464 <= 0;
      __delay_data_2022_greaterthan_1460 <= 0;
      __delay_data_2023_greatereq_1473 <= 0;
      __delay_data_2026__delay_2025__variable_1457 <= 0;
      __delay_data_2029__delay_2028__variable_1458 <= 0;
      __delay_data_2032__delay_2031__variable_1459 <= 0;
      _cond_data_1470 <= 0;
      __delay_data_2024__delay_2023_greatereq_1473 <= 0;
      __delay_data_2027__delay_2026__delay_2025__variable_1457 <= 0;
      __delay_data_2030__delay_2029__delay_2028__variable_1458 <= 0;
      __delay_data_2033__delay_2032__delay_2031__variable_1459 <= 0;
      __muladd_madd_odata_reg_1476 <= 0;
      __delay_data_2034__delay_2033__delay_2032____variable_1459 <= 0;
      __delay_data_2035__delay_2034__delay_2033____variable_1459 <= 0;
      __delay_data_2036__delay_2035__delay_2034____variable_1459 <= 0;
      __delay_data_2037__delay_2036__delay_2035____variable_1459 <= 0;
      _sra_data_1477 <= 0;
      __variable_wdata_1457 <= 0;
      __variable_wdata_1458 <= 0;
      __variable_wdata_1459 <= 0;
      _tmp_799 <= 0;
      _tmp_800 <= 0;
      _tmp_801 <= 0;
      _tmp_802 <= 0;
      _tmp_803 <= 0;
      _tmp_804 <= 0;
      _tmp_805 <= 0;
      _tmp_806 <= 0;
      _tmp_807 <= 0;
      _tmp_808 <= 0;
      _tmp_809 <= 0;
      _tmp_810 <= 0;
      _tmp_811 <= 0;
      _tmp_812 <= 0;
      _tmp_813 <= 0;
      _tmp_814 <= 0;
      _tmp_815 <= 0;
      _tmp_816 <= 0;
      _tmp_817 <= 0;
      _tmp_818 <= 0;
      _tmp_819 <= 0;
      _tmp_820 <= 0;
      _tmp_821 <= 0;
      _tmp_822 <= 0;
      _tmp_823 <= 0;
      _tmp_824 <= 0;
      _tmp_825 <= 0;
      _tmp_826 <= 0;
      _tmp_827 <= 0;
      _tmp_828 <= 0;
      _tmp_829 <= 0;
      _tmp_830 <= 0;
      _tmp_831 <= 0;
      _tmp_832 <= 0;
      _mul_23_busy_reg <= 0;
    end else begin
      if(_mul_23_stream_oready) begin
        _mul_23_x_source_ram_renable <= 0;
        _mul_23_x_source_fifo_deq <= 0;
      end 
      _mul_23_x_idle <= _mul_23_x_idle;
      if(_mul_23_stream_oready) begin
        _mul_23_y_source_ram_renable <= 0;
        _mul_23_y_source_fifo_deq <= 0;
      end 
      _mul_23_y_idle <= _mul_23_y_idle;
      if(_mul_23_stream_oready) begin
        _mul_23_rshift_source_ram_renable <= 0;
        _mul_23_rshift_source_fifo_deq <= 0;
      end 
      _mul_23_rshift_idle <= _mul_23_rshift_idle;
      if(_mul_23_stream_oready) begin
        _mul_23_z_sink_wenable <= 0;
        _mul_23_z_sink_fifo_enq <= 0;
      end 
      if(_mul_23_stream_oready) begin
        __mul_23_stream_ivalid_1 <= _mul_23_stream_ivalid;
      end 
      if(_mul_23_stream_oready) begin
        __mul_23_stream_ivalid_2 <= __mul_23_stream_ivalid_1;
      end 
      if(_mul_23_stream_oready) begin
        __mul_23_stream_ivalid_3 <= __mul_23_stream_ivalid_2;
      end 
      if(_mul_23_stream_oready) begin
        __mul_23_stream_ivalid_4 <= __mul_23_stream_ivalid_3;
      end 
      if(_mul_23_stream_oready) begin
        __mul_23_stream_ivalid_5 <= __mul_23_stream_ivalid_4;
      end 
      if(_mul_23_stream_oready) begin
        __mul_23_stream_ivalid_6 <= __mul_23_stream_ivalid_5;
      end 
      if(_mul_23_stream_oready) begin
        __mul_23_stream_ivalid_7 <= __mul_23_stream_ivalid_6;
      end 
      if(_mul_23_stream_oready) begin
        __mul_23_stream_ivalid_8 <= __mul_23_stream_ivalid_7;
      end 
      if(_mul_23_stream_oready) begin
        _greaterthan_data_1460 <= mul_23_rshift_data > 1'sd0;
      end 
      if(_mul_23_stream_oready) begin
        _minus_data_1462 <= mul_23_rshift_data - 2'sd1;
      end 
      if(_mul_23_stream_oready) begin
        _greatereq_data_1473 <= mul_23_x_data >= 1'sd0;
      end 
      if(_mul_23_stream_oready) begin
        __delay_data_2025__variable_1457 <= mul_23_x_data;
      end 
      if(_mul_23_stream_oready) begin
        __delay_data_2028__variable_1458 <= mul_23_y_data;
      end 
      if(_mul_23_stream_oready) begin
        __delay_data_2031__variable_1459 <= mul_23_rshift_data;
      end 
      if(_mul_23_stream_oready) begin
        _sll_data_1464 <= 2'sd1 << _minus_data_1462;
      end 
      if(_mul_23_stream_oready) begin
        __delay_data_2022_greaterthan_1460 <= _greaterthan_data_1460;
      end 
      if(_mul_23_stream_oready) begin
        __delay_data_2023_greatereq_1473 <= _greatereq_data_1473;
      end 
      if(_mul_23_stream_oready) begin
        __delay_data_2026__delay_2025__variable_1457 <= __delay_data_2025__variable_1457;
      end 
      if(_mul_23_stream_oready) begin
        __delay_data_2029__delay_2028__variable_1458 <= __delay_data_2028__variable_1458;
      end 
      if(_mul_23_stream_oready) begin
        __delay_data_2032__delay_2031__variable_1459 <= __delay_data_2031__variable_1459;
      end 
      if(_mul_23_stream_oready) begin
        _cond_data_1470 <= (__delay_data_2022_greaterthan_1460)? _sll_data_1464 : 1'sd0;
      end 
      if(_mul_23_stream_oready) begin
        __delay_data_2024__delay_2023_greatereq_1473 <= __delay_data_2023_greatereq_1473;
      end 
      if(_mul_23_stream_oready) begin
        __delay_data_2027__delay_2026__delay_2025__variable_1457 <= __delay_data_2026__delay_2025__variable_1457;
      end 
      if(_mul_23_stream_oready) begin
        __delay_data_2030__delay_2029__delay_2028__variable_1458 <= __delay_data_2029__delay_2028__variable_1458;
      end 
      if(_mul_23_stream_oready) begin
        __delay_data_2033__delay_2032__delay_2031__variable_1459 <= __delay_data_2032__delay_2031__variable_1459;
      end 
      if(_mul_23_stream_oready) begin
        __muladd_madd_odata_reg_1476 <= __muladd_madd_odata_1476;
      end 
      if(_mul_23_stream_oready) begin
        __delay_data_2034__delay_2033__delay_2032____variable_1459 <= __delay_data_2033__delay_2032__delay_2031__variable_1459;
      end 
      if(_mul_23_stream_oready) begin
        __delay_data_2035__delay_2034__delay_2033____variable_1459 <= __delay_data_2034__delay_2033__delay_2032____variable_1459;
      end 
      if(_mul_23_stream_oready) begin
        __delay_data_2036__delay_2035__delay_2034____variable_1459 <= __delay_data_2035__delay_2034__delay_2033____variable_1459;
      end 
      if(_mul_23_stream_oready) begin
        __delay_data_2037__delay_2036__delay_2035____variable_1459 <= __delay_data_2036__delay_2035__delay_2034____variable_1459;
      end 
      if(_mul_23_stream_oready) begin
        _sra_data_1477 <= __muladd_data_1476 >>> __delay_data_2037__delay_2036__delay_2035____variable_1459;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_1457 <= _cond_data_1919;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_1458 <= __delay_data_2278_reinterpretcast_1886;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_1459 <= _plus_data_2038;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_799 <= _mul_23_source_start;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_800 <= _tmp_799;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_801 <= _tmp_800;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_802 <= _mul_23_source_start;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_803 <= _tmp_802;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_804 <= _tmp_803;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_805 <= _tmp_804;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_806 <= _tmp_805;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_807 <= _tmp_806;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_808 <= _tmp_807;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_809 <= _tmp_808;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_810 <= _tmp_809;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_811 <= _tmp_810;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_812 <= _mul_23_source_stop;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_813 <= _tmp_812;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_814 <= _tmp_813;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_815 <= _tmp_814;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_816 <= _tmp_815;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_817 <= _tmp_816;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_818 <= _tmp_817;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_819 <= _tmp_818;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_820 <= _tmp_819;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_821 <= _tmp_820;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_822 <= _mul_23_source_busy;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_823 <= _tmp_822;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_824 <= _tmp_823;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_825 <= _tmp_824;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_826 <= _tmp_825;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_827 <= _tmp_826;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_828 <= _tmp_827;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_829 <= _tmp_828;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_830 <= _tmp_829;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_831 <= _tmp_830;
      end 
      if(_mul_23_stream_oready) begin
        _tmp_832 <= _mul_23_sink_busy;
      end 
      if(!_mul_23_sink_busy && _tmp_832) begin
        _mul_23_busy_reg <= 0;
      end 
      if(_mul_23_source_busy) begin
        _mul_23_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_23_fsm_1 = 1;
  localparam _mul_23_fsm_2 = 2;
  localparam _mul_23_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_23_fsm <= _mul_23_fsm_init;
      _mul_23_source_start <= 0;
      _mul_23_source_busy <= 0;
      _mul_23_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        _mul_23_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_23_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_23_stream_oready && _tmp_801) begin
        _mul_23_stream_ivalid <= 1;
      end 
      if(_mul_23_stream_oready && 1'd0) begin
        _mul_23_stream_ivalid <= 0;
      end 
      case(_mul_23_fsm)
        _mul_23_fsm_init: begin
          if(_mul_23_run_flag) begin
            _mul_23_source_start <= 1;
          end 
          if(_mul_23_run_flag) begin
            _mul_23_fsm <= _mul_23_fsm_1;
          end 
        end
        _mul_23_fsm_1: begin
          if(_mul_23_source_start && _mul_23_stream_oready) begin
            _mul_23_source_start <= 0;
            _mul_23_source_busy <= 1;
          end 
          if(_mul_23_source_start && _mul_23_stream_oready) begin
            _mul_23_fsm <= _mul_23_fsm_2;
          end 
        end
        _mul_23_fsm_2: begin
          if(_mul_23_stream_oready) begin
            _mul_23_fsm <= _mul_23_fsm_3;
          end 
        end
        _mul_23_fsm_3: begin
          if(_mul_23_stream_oready && 1'd0) begin
            _mul_23_source_busy <= 0;
          end 
          if(_mul_23_stream_oready && 1'd0 && _mul_23_run_flag) begin
            _mul_23_source_start <= 1;
          end 
          if(_mul_23_stream_oready && 1'd0) begin
            _mul_23_fsm <= _mul_23_fsm_init;
          end 
          if(_mul_23_stream_oready && 1'd0 && _mul_23_run_flag) begin
            _mul_23_fsm <= _mul_23_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_24_x_source_ram_renable <= 0;
      _mul_24_x_source_fifo_deq <= 0;
      _mul_24_x_idle <= 1;
      _mul_24_y_source_ram_renable <= 0;
      _mul_24_y_source_fifo_deq <= 0;
      _mul_24_y_idle <= 1;
      _mul_24_rshift_source_ram_renable <= 0;
      _mul_24_rshift_source_fifo_deq <= 0;
      _mul_24_rshift_idle <= 1;
      _mul_24_z_sink_wenable <= 0;
      _mul_24_z_sink_fifo_enq <= 0;
      __mul_24_stream_ivalid_1 <= 0;
      __mul_24_stream_ivalid_2 <= 0;
      __mul_24_stream_ivalid_3 <= 0;
      __mul_24_stream_ivalid_4 <= 0;
      __mul_24_stream_ivalid_5 <= 0;
      __mul_24_stream_ivalid_6 <= 0;
      __mul_24_stream_ivalid_7 <= 0;
      __mul_24_stream_ivalid_8 <= 0;
      _greaterthan_data_1481 <= 0;
      _minus_data_1483 <= 0;
      _greatereq_data_1494 <= 0;
      __delay_data_2044__variable_1478 <= 0;
      __delay_data_2047__variable_1479 <= 0;
      __delay_data_2050__variable_1480 <= 0;
      _sll_data_1485 <= 0;
      __delay_data_2041_greaterthan_1481 <= 0;
      __delay_data_2042_greatereq_1494 <= 0;
      __delay_data_2045__delay_2044__variable_1478 <= 0;
      __delay_data_2048__delay_2047__variable_1479 <= 0;
      __delay_data_2051__delay_2050__variable_1480 <= 0;
      _cond_data_1491 <= 0;
      __delay_data_2043__delay_2042_greatereq_1494 <= 0;
      __delay_data_2046__delay_2045__delay_2044__variable_1478 <= 0;
      __delay_data_2049__delay_2048__delay_2047__variable_1479 <= 0;
      __delay_data_2052__delay_2051__delay_2050__variable_1480 <= 0;
      __muladd_madd_odata_reg_1497 <= 0;
      __delay_data_2053__delay_2052__delay_2051____variable_1480 <= 0;
      __delay_data_2054__delay_2053__delay_2052____variable_1480 <= 0;
      __delay_data_2055__delay_2054__delay_2053____variable_1480 <= 0;
      __delay_data_2056__delay_2055__delay_2054____variable_1480 <= 0;
      _sra_data_1498 <= 0;
      __variable_wdata_1478 <= 0;
      __variable_wdata_1479 <= 0;
      __variable_wdata_1480 <= 0;
      _tmp_833 <= 0;
      _tmp_834 <= 0;
      _tmp_835 <= 0;
      _tmp_836 <= 0;
      _tmp_837 <= 0;
      _tmp_838 <= 0;
      _tmp_839 <= 0;
      _tmp_840 <= 0;
      _tmp_841 <= 0;
      _tmp_842 <= 0;
      _tmp_843 <= 0;
      _tmp_844 <= 0;
      _tmp_845 <= 0;
      _tmp_846 <= 0;
      _tmp_847 <= 0;
      _tmp_848 <= 0;
      _tmp_849 <= 0;
      _tmp_850 <= 0;
      _tmp_851 <= 0;
      _tmp_852 <= 0;
      _tmp_853 <= 0;
      _tmp_854 <= 0;
      _tmp_855 <= 0;
      _tmp_856 <= 0;
      _tmp_857 <= 0;
      _tmp_858 <= 0;
      _tmp_859 <= 0;
      _tmp_860 <= 0;
      _tmp_861 <= 0;
      _tmp_862 <= 0;
      _tmp_863 <= 0;
      _tmp_864 <= 0;
      _tmp_865 <= 0;
      _tmp_866 <= 0;
      _mul_24_busy_reg <= 0;
    end else begin
      if(_mul_24_stream_oready) begin
        _mul_24_x_source_ram_renable <= 0;
        _mul_24_x_source_fifo_deq <= 0;
      end 
      _mul_24_x_idle <= _mul_24_x_idle;
      if(_mul_24_stream_oready) begin
        _mul_24_y_source_ram_renable <= 0;
        _mul_24_y_source_fifo_deq <= 0;
      end 
      _mul_24_y_idle <= _mul_24_y_idle;
      if(_mul_24_stream_oready) begin
        _mul_24_rshift_source_ram_renable <= 0;
        _mul_24_rshift_source_fifo_deq <= 0;
      end 
      _mul_24_rshift_idle <= _mul_24_rshift_idle;
      if(_mul_24_stream_oready) begin
        _mul_24_z_sink_wenable <= 0;
        _mul_24_z_sink_fifo_enq <= 0;
      end 
      if(_mul_24_stream_oready) begin
        __mul_24_stream_ivalid_1 <= _mul_24_stream_ivalid;
      end 
      if(_mul_24_stream_oready) begin
        __mul_24_stream_ivalid_2 <= __mul_24_stream_ivalid_1;
      end 
      if(_mul_24_stream_oready) begin
        __mul_24_stream_ivalid_3 <= __mul_24_stream_ivalid_2;
      end 
      if(_mul_24_stream_oready) begin
        __mul_24_stream_ivalid_4 <= __mul_24_stream_ivalid_3;
      end 
      if(_mul_24_stream_oready) begin
        __mul_24_stream_ivalid_5 <= __mul_24_stream_ivalid_4;
      end 
      if(_mul_24_stream_oready) begin
        __mul_24_stream_ivalid_6 <= __mul_24_stream_ivalid_5;
      end 
      if(_mul_24_stream_oready) begin
        __mul_24_stream_ivalid_7 <= __mul_24_stream_ivalid_6;
      end 
      if(_mul_24_stream_oready) begin
        __mul_24_stream_ivalid_8 <= __mul_24_stream_ivalid_7;
      end 
      if(_mul_24_stream_oready) begin
        _greaterthan_data_1481 <= mul_24_rshift_data > 1'sd0;
      end 
      if(_mul_24_stream_oready) begin
        _minus_data_1483 <= mul_24_rshift_data - 2'sd1;
      end 
      if(_mul_24_stream_oready) begin
        _greatereq_data_1494 <= mul_24_x_data >= 1'sd0;
      end 
      if(_mul_24_stream_oready) begin
        __delay_data_2044__variable_1478 <= mul_24_x_data;
      end 
      if(_mul_24_stream_oready) begin
        __delay_data_2047__variable_1479 <= mul_24_y_data;
      end 
      if(_mul_24_stream_oready) begin
        __delay_data_2050__variable_1480 <= mul_24_rshift_data;
      end 
      if(_mul_24_stream_oready) begin
        _sll_data_1485 <= 2'sd1 << _minus_data_1483;
      end 
      if(_mul_24_stream_oready) begin
        __delay_data_2041_greaterthan_1481 <= _greaterthan_data_1481;
      end 
      if(_mul_24_stream_oready) begin
        __delay_data_2042_greatereq_1494 <= _greatereq_data_1494;
      end 
      if(_mul_24_stream_oready) begin
        __delay_data_2045__delay_2044__variable_1478 <= __delay_data_2044__variable_1478;
      end 
      if(_mul_24_stream_oready) begin
        __delay_data_2048__delay_2047__variable_1479 <= __delay_data_2047__variable_1479;
      end 
      if(_mul_24_stream_oready) begin
        __delay_data_2051__delay_2050__variable_1480 <= __delay_data_2050__variable_1480;
      end 
      if(_mul_24_stream_oready) begin
        _cond_data_1491 <= (__delay_data_2041_greaterthan_1481)? _sll_data_1485 : 1'sd0;
      end 
      if(_mul_24_stream_oready) begin
        __delay_data_2043__delay_2042_greatereq_1494 <= __delay_data_2042_greatereq_1494;
      end 
      if(_mul_24_stream_oready) begin
        __delay_data_2046__delay_2045__delay_2044__variable_1478 <= __delay_data_2045__delay_2044__variable_1478;
      end 
      if(_mul_24_stream_oready) begin
        __delay_data_2049__delay_2048__delay_2047__variable_1479 <= __delay_data_2048__delay_2047__variable_1479;
      end 
      if(_mul_24_stream_oready) begin
        __delay_data_2052__delay_2051__delay_2050__variable_1480 <= __delay_data_2051__delay_2050__variable_1480;
      end 
      if(_mul_24_stream_oready) begin
        __muladd_madd_odata_reg_1497 <= __muladd_madd_odata_1497;
      end 
      if(_mul_24_stream_oready) begin
        __delay_data_2053__delay_2052__delay_2051____variable_1480 <= __delay_data_2052__delay_2051__delay_2050__variable_1480;
      end 
      if(_mul_24_stream_oready) begin
        __delay_data_2054__delay_2053__delay_2052____variable_1480 <= __delay_data_2053__delay_2052__delay_2051____variable_1480;
      end 
      if(_mul_24_stream_oready) begin
        __delay_data_2055__delay_2054__delay_2053____variable_1480 <= __delay_data_2054__delay_2053__delay_2052____variable_1480;
      end 
      if(_mul_24_stream_oready) begin
        __delay_data_2056__delay_2055__delay_2054____variable_1480 <= __delay_data_2055__delay_2054__delay_2053____variable_1480;
      end 
      if(_mul_24_stream_oready) begin
        _sra_data_1498 <= __muladd_data_1497 >>> __delay_data_2056__delay_2055__delay_2054____variable_1480;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_1478 <= _cond_data_1921;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_1479 <= __delay_data_2280_reinterpretcast_1887;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_1480 <= _plus_data_2057;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_833 <= _mul_24_source_start;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_834 <= _tmp_833;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_835 <= _tmp_834;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_836 <= _mul_24_source_start;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_837 <= _tmp_836;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_838 <= _tmp_837;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_839 <= _tmp_838;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_840 <= _tmp_839;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_841 <= _tmp_840;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_842 <= _tmp_841;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_843 <= _tmp_842;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_844 <= _tmp_843;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_845 <= _tmp_844;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_846 <= _mul_24_source_stop;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_847 <= _tmp_846;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_848 <= _tmp_847;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_849 <= _tmp_848;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_850 <= _tmp_849;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_851 <= _tmp_850;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_852 <= _tmp_851;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_853 <= _tmp_852;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_854 <= _tmp_853;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_855 <= _tmp_854;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_856 <= _mul_24_source_busy;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_857 <= _tmp_856;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_858 <= _tmp_857;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_859 <= _tmp_858;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_860 <= _tmp_859;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_861 <= _tmp_860;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_862 <= _tmp_861;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_863 <= _tmp_862;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_864 <= _tmp_863;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_865 <= _tmp_864;
      end 
      if(_mul_24_stream_oready) begin
        _tmp_866 <= _mul_24_sink_busy;
      end 
      if(!_mul_24_sink_busy && _tmp_866) begin
        _mul_24_busy_reg <= 0;
      end 
      if(_mul_24_source_busy) begin
        _mul_24_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_24_fsm_1 = 1;
  localparam _mul_24_fsm_2 = 2;
  localparam _mul_24_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_24_fsm <= _mul_24_fsm_init;
      _mul_24_source_start <= 0;
      _mul_24_source_busy <= 0;
      _mul_24_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        _mul_24_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_24_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_24_stream_oready && _tmp_835) begin
        _mul_24_stream_ivalid <= 1;
      end 
      if(_mul_24_stream_oready && 1'd0) begin
        _mul_24_stream_ivalid <= 0;
      end 
      case(_mul_24_fsm)
        _mul_24_fsm_init: begin
          if(_mul_24_run_flag) begin
            _mul_24_source_start <= 1;
          end 
          if(_mul_24_run_flag) begin
            _mul_24_fsm <= _mul_24_fsm_1;
          end 
        end
        _mul_24_fsm_1: begin
          if(_mul_24_source_start && _mul_24_stream_oready) begin
            _mul_24_source_start <= 0;
            _mul_24_source_busy <= 1;
          end 
          if(_mul_24_source_start && _mul_24_stream_oready) begin
            _mul_24_fsm <= _mul_24_fsm_2;
          end 
        end
        _mul_24_fsm_2: begin
          if(_mul_24_stream_oready) begin
            _mul_24_fsm <= _mul_24_fsm_3;
          end 
        end
        _mul_24_fsm_3: begin
          if(_mul_24_stream_oready && 1'd0) begin
            _mul_24_source_busy <= 0;
          end 
          if(_mul_24_stream_oready && 1'd0 && _mul_24_run_flag) begin
            _mul_24_source_start <= 1;
          end 
          if(_mul_24_stream_oready && 1'd0) begin
            _mul_24_fsm <= _mul_24_fsm_init;
          end 
          if(_mul_24_stream_oready && 1'd0 && _mul_24_run_flag) begin
            _mul_24_fsm <= _mul_24_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_25_x_source_ram_renable <= 0;
      _mul_25_x_source_fifo_deq <= 0;
      _mul_25_x_idle <= 1;
      _mul_25_y_source_ram_renable <= 0;
      _mul_25_y_source_fifo_deq <= 0;
      _mul_25_y_idle <= 1;
      _mul_25_rshift_source_ram_renable <= 0;
      _mul_25_rshift_source_fifo_deq <= 0;
      _mul_25_rshift_idle <= 1;
      _mul_25_z_sink_wenable <= 0;
      _mul_25_z_sink_fifo_enq <= 0;
      __mul_25_stream_ivalid_1 <= 0;
      __mul_25_stream_ivalid_2 <= 0;
      __mul_25_stream_ivalid_3 <= 0;
      __mul_25_stream_ivalid_4 <= 0;
      __mul_25_stream_ivalid_5 <= 0;
      __mul_25_stream_ivalid_6 <= 0;
      __mul_25_stream_ivalid_7 <= 0;
      __mul_25_stream_ivalid_8 <= 0;
      _greaterthan_data_1502 <= 0;
      _minus_data_1504 <= 0;
      _greatereq_data_1515 <= 0;
      __delay_data_2063__variable_1499 <= 0;
      __delay_data_2066__variable_1500 <= 0;
      __delay_data_2069__variable_1501 <= 0;
      _sll_data_1506 <= 0;
      __delay_data_2060_greaterthan_1502 <= 0;
      __delay_data_2061_greatereq_1515 <= 0;
      __delay_data_2064__delay_2063__variable_1499 <= 0;
      __delay_data_2067__delay_2066__variable_1500 <= 0;
      __delay_data_2070__delay_2069__variable_1501 <= 0;
      _cond_data_1512 <= 0;
      __delay_data_2062__delay_2061_greatereq_1515 <= 0;
      __delay_data_2065__delay_2064__delay_2063__variable_1499 <= 0;
      __delay_data_2068__delay_2067__delay_2066__variable_1500 <= 0;
      __delay_data_2071__delay_2070__delay_2069__variable_1501 <= 0;
      __muladd_madd_odata_reg_1518 <= 0;
      __delay_data_2072__delay_2071__delay_2070____variable_1501 <= 0;
      __delay_data_2073__delay_2072__delay_2071____variable_1501 <= 0;
      __delay_data_2074__delay_2073__delay_2072____variable_1501 <= 0;
      __delay_data_2075__delay_2074__delay_2073____variable_1501 <= 0;
      _sra_data_1519 <= 0;
      __variable_wdata_1499 <= 0;
      __variable_wdata_1500 <= 0;
      __variable_wdata_1501 <= 0;
      _tmp_867 <= 0;
      _tmp_868 <= 0;
      _tmp_869 <= 0;
      _tmp_870 <= 0;
      _tmp_871 <= 0;
      _tmp_872 <= 0;
      _tmp_873 <= 0;
      _tmp_874 <= 0;
      _tmp_875 <= 0;
      _tmp_876 <= 0;
      _tmp_877 <= 0;
      _tmp_878 <= 0;
      _tmp_879 <= 0;
      _tmp_880 <= 0;
      _tmp_881 <= 0;
      _tmp_882 <= 0;
      _tmp_883 <= 0;
      _tmp_884 <= 0;
      _tmp_885 <= 0;
      _tmp_886 <= 0;
      _tmp_887 <= 0;
      _tmp_888 <= 0;
      _tmp_889 <= 0;
      _tmp_890 <= 0;
      _tmp_891 <= 0;
      _tmp_892 <= 0;
      _tmp_893 <= 0;
      _tmp_894 <= 0;
      _tmp_895 <= 0;
      _tmp_896 <= 0;
      _tmp_897 <= 0;
      _tmp_898 <= 0;
      _tmp_899 <= 0;
      _tmp_900 <= 0;
      _mul_25_busy_reg <= 0;
    end else begin
      if(_mul_25_stream_oready) begin
        _mul_25_x_source_ram_renable <= 0;
        _mul_25_x_source_fifo_deq <= 0;
      end 
      _mul_25_x_idle <= _mul_25_x_idle;
      if(_mul_25_stream_oready) begin
        _mul_25_y_source_ram_renable <= 0;
        _mul_25_y_source_fifo_deq <= 0;
      end 
      _mul_25_y_idle <= _mul_25_y_idle;
      if(_mul_25_stream_oready) begin
        _mul_25_rshift_source_ram_renable <= 0;
        _mul_25_rshift_source_fifo_deq <= 0;
      end 
      _mul_25_rshift_idle <= _mul_25_rshift_idle;
      if(_mul_25_stream_oready) begin
        _mul_25_z_sink_wenable <= 0;
        _mul_25_z_sink_fifo_enq <= 0;
      end 
      if(_mul_25_stream_oready) begin
        __mul_25_stream_ivalid_1 <= _mul_25_stream_ivalid;
      end 
      if(_mul_25_stream_oready) begin
        __mul_25_stream_ivalid_2 <= __mul_25_stream_ivalid_1;
      end 
      if(_mul_25_stream_oready) begin
        __mul_25_stream_ivalid_3 <= __mul_25_stream_ivalid_2;
      end 
      if(_mul_25_stream_oready) begin
        __mul_25_stream_ivalid_4 <= __mul_25_stream_ivalid_3;
      end 
      if(_mul_25_stream_oready) begin
        __mul_25_stream_ivalid_5 <= __mul_25_stream_ivalid_4;
      end 
      if(_mul_25_stream_oready) begin
        __mul_25_stream_ivalid_6 <= __mul_25_stream_ivalid_5;
      end 
      if(_mul_25_stream_oready) begin
        __mul_25_stream_ivalid_7 <= __mul_25_stream_ivalid_6;
      end 
      if(_mul_25_stream_oready) begin
        __mul_25_stream_ivalid_8 <= __mul_25_stream_ivalid_7;
      end 
      if(_mul_25_stream_oready) begin
        _greaterthan_data_1502 <= mul_25_rshift_data > 1'sd0;
      end 
      if(_mul_25_stream_oready) begin
        _minus_data_1504 <= mul_25_rshift_data - 2'sd1;
      end 
      if(_mul_25_stream_oready) begin
        _greatereq_data_1515 <= mul_25_x_data >= 1'sd0;
      end 
      if(_mul_25_stream_oready) begin
        __delay_data_2063__variable_1499 <= mul_25_x_data;
      end 
      if(_mul_25_stream_oready) begin
        __delay_data_2066__variable_1500 <= mul_25_y_data;
      end 
      if(_mul_25_stream_oready) begin
        __delay_data_2069__variable_1501 <= mul_25_rshift_data;
      end 
      if(_mul_25_stream_oready) begin
        _sll_data_1506 <= 2'sd1 << _minus_data_1504;
      end 
      if(_mul_25_stream_oready) begin
        __delay_data_2060_greaterthan_1502 <= _greaterthan_data_1502;
      end 
      if(_mul_25_stream_oready) begin
        __delay_data_2061_greatereq_1515 <= _greatereq_data_1515;
      end 
      if(_mul_25_stream_oready) begin
        __delay_data_2064__delay_2063__variable_1499 <= __delay_data_2063__variable_1499;
      end 
      if(_mul_25_stream_oready) begin
        __delay_data_2067__delay_2066__variable_1500 <= __delay_data_2066__variable_1500;
      end 
      if(_mul_25_stream_oready) begin
        __delay_data_2070__delay_2069__variable_1501 <= __delay_data_2069__variable_1501;
      end 
      if(_mul_25_stream_oready) begin
        _cond_data_1512 <= (__delay_data_2060_greaterthan_1502)? _sll_data_1506 : 1'sd0;
      end 
      if(_mul_25_stream_oready) begin
        __delay_data_2062__delay_2061_greatereq_1515 <= __delay_data_2061_greatereq_1515;
      end 
      if(_mul_25_stream_oready) begin
        __delay_data_2065__delay_2064__delay_2063__variable_1499 <= __delay_data_2064__delay_2063__variable_1499;
      end 
      if(_mul_25_stream_oready) begin
        __delay_data_2068__delay_2067__delay_2066__variable_1500 <= __delay_data_2067__delay_2066__variable_1500;
      end 
      if(_mul_25_stream_oready) begin
        __delay_data_2071__delay_2070__delay_2069__variable_1501 <= __delay_data_2070__delay_2069__variable_1501;
      end 
      if(_mul_25_stream_oready) begin
        __muladd_madd_odata_reg_1518 <= __muladd_madd_odata_1518;
      end 
      if(_mul_25_stream_oready) begin
        __delay_data_2072__delay_2071__delay_2070____variable_1501 <= __delay_data_2071__delay_2070__delay_2069__variable_1501;
      end 
      if(_mul_25_stream_oready) begin
        __delay_data_2073__delay_2072__delay_2071____variable_1501 <= __delay_data_2072__delay_2071__delay_2070____variable_1501;
      end 
      if(_mul_25_stream_oready) begin
        __delay_data_2074__delay_2073__delay_2072____variable_1501 <= __delay_data_2073__delay_2072__delay_2071____variable_1501;
      end 
      if(_mul_25_stream_oready) begin
        __delay_data_2075__delay_2074__delay_2073____variable_1501 <= __delay_data_2074__delay_2073__delay_2072____variable_1501;
      end 
      if(_mul_25_stream_oready) begin
        _sra_data_1519 <= __muladd_data_1518 >>> __delay_data_2075__delay_2074__delay_2073____variable_1501;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_1499 <= _cond_data_1923;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_1500 <= __delay_data_2282_reinterpretcast_1888;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_1501 <= _plus_data_2076;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_867 <= _mul_25_source_start;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_868 <= _tmp_867;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_869 <= _tmp_868;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_870 <= _mul_25_source_start;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_871 <= _tmp_870;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_872 <= _tmp_871;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_873 <= _tmp_872;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_874 <= _tmp_873;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_875 <= _tmp_874;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_876 <= _tmp_875;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_877 <= _tmp_876;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_878 <= _tmp_877;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_879 <= _tmp_878;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_880 <= _mul_25_source_stop;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_881 <= _tmp_880;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_882 <= _tmp_881;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_883 <= _tmp_882;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_884 <= _tmp_883;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_885 <= _tmp_884;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_886 <= _tmp_885;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_887 <= _tmp_886;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_888 <= _tmp_887;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_889 <= _tmp_888;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_890 <= _mul_25_source_busy;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_891 <= _tmp_890;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_892 <= _tmp_891;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_893 <= _tmp_892;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_894 <= _tmp_893;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_895 <= _tmp_894;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_896 <= _tmp_895;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_897 <= _tmp_896;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_898 <= _tmp_897;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_899 <= _tmp_898;
      end 
      if(_mul_25_stream_oready) begin
        _tmp_900 <= _mul_25_sink_busy;
      end 
      if(!_mul_25_sink_busy && _tmp_900) begin
        _mul_25_busy_reg <= 0;
      end 
      if(_mul_25_source_busy) begin
        _mul_25_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_25_fsm_1 = 1;
  localparam _mul_25_fsm_2 = 2;
  localparam _mul_25_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_25_fsm <= _mul_25_fsm_init;
      _mul_25_source_start <= 0;
      _mul_25_source_busy <= 0;
      _mul_25_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        _mul_25_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_25_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_25_stream_oready && _tmp_869) begin
        _mul_25_stream_ivalid <= 1;
      end 
      if(_mul_25_stream_oready && 1'd0) begin
        _mul_25_stream_ivalid <= 0;
      end 
      case(_mul_25_fsm)
        _mul_25_fsm_init: begin
          if(_mul_25_run_flag) begin
            _mul_25_source_start <= 1;
          end 
          if(_mul_25_run_flag) begin
            _mul_25_fsm <= _mul_25_fsm_1;
          end 
        end
        _mul_25_fsm_1: begin
          if(_mul_25_source_start && _mul_25_stream_oready) begin
            _mul_25_source_start <= 0;
            _mul_25_source_busy <= 1;
          end 
          if(_mul_25_source_start && _mul_25_stream_oready) begin
            _mul_25_fsm <= _mul_25_fsm_2;
          end 
        end
        _mul_25_fsm_2: begin
          if(_mul_25_stream_oready) begin
            _mul_25_fsm <= _mul_25_fsm_3;
          end 
        end
        _mul_25_fsm_3: begin
          if(_mul_25_stream_oready && 1'd0) begin
            _mul_25_source_busy <= 0;
          end 
          if(_mul_25_stream_oready && 1'd0 && _mul_25_run_flag) begin
            _mul_25_source_start <= 1;
          end 
          if(_mul_25_stream_oready && 1'd0) begin
            _mul_25_fsm <= _mul_25_fsm_init;
          end 
          if(_mul_25_stream_oready && 1'd0 && _mul_25_run_flag) begin
            _mul_25_fsm <= _mul_25_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mul_26_x_source_ram_renable <= 0;
      _mul_26_x_source_fifo_deq <= 0;
      _mul_26_x_idle <= 1;
      _mul_26_y_source_ram_renable <= 0;
      _mul_26_y_source_fifo_deq <= 0;
      _mul_26_y_idle <= 1;
      _mul_26_rshift_source_ram_renable <= 0;
      _mul_26_rshift_source_fifo_deq <= 0;
      _mul_26_rshift_idle <= 1;
      _mul_26_z_sink_wenable <= 0;
      _mul_26_z_sink_fifo_enq <= 0;
      __mul_26_stream_ivalid_1 <= 0;
      __mul_26_stream_ivalid_2 <= 0;
      __mul_26_stream_ivalid_3 <= 0;
      __mul_26_stream_ivalid_4 <= 0;
      __mul_26_stream_ivalid_5 <= 0;
      __mul_26_stream_ivalid_6 <= 0;
      __mul_26_stream_ivalid_7 <= 0;
      __mul_26_stream_ivalid_8 <= 0;
      _greaterthan_data_1523 <= 0;
      _minus_data_1525 <= 0;
      _greatereq_data_1536 <= 0;
      __delay_data_2082__variable_1520 <= 0;
      __delay_data_2085__variable_1521 <= 0;
      __delay_data_2088__variable_1522 <= 0;
      _sll_data_1527 <= 0;
      __delay_data_2079_greaterthan_1523 <= 0;
      __delay_data_2080_greatereq_1536 <= 0;
      __delay_data_2083__delay_2082__variable_1520 <= 0;
      __delay_data_2086__delay_2085__variable_1521 <= 0;
      __delay_data_2089__delay_2088__variable_1522 <= 0;
      _cond_data_1533 <= 0;
      __delay_data_2081__delay_2080_greatereq_1536 <= 0;
      __delay_data_2084__delay_2083__delay_2082__variable_1520 <= 0;
      __delay_data_2087__delay_2086__delay_2085__variable_1521 <= 0;
      __delay_data_2090__delay_2089__delay_2088__variable_1522 <= 0;
      __muladd_madd_odata_reg_1539 <= 0;
      __delay_data_2091__delay_2090__delay_2089____variable_1522 <= 0;
      __delay_data_2092__delay_2091__delay_2090____variable_1522 <= 0;
      __delay_data_2093__delay_2092__delay_2091____variable_1522 <= 0;
      __delay_data_2094__delay_2093__delay_2092____variable_1522 <= 0;
      _sra_data_1540 <= 0;
      __variable_wdata_1520 <= 0;
      __variable_wdata_1521 <= 0;
      __variable_wdata_1522 <= 0;
      _tmp_901 <= 0;
      _tmp_902 <= 0;
      _tmp_903 <= 0;
      _tmp_904 <= 0;
      _tmp_905 <= 0;
      _tmp_906 <= 0;
      _tmp_907 <= 0;
      _tmp_908 <= 0;
      _tmp_909 <= 0;
      _tmp_910 <= 0;
      _tmp_911 <= 0;
      _tmp_912 <= 0;
      _tmp_913 <= 0;
      _tmp_914 <= 0;
      _tmp_915 <= 0;
      _tmp_916 <= 0;
      _tmp_917 <= 0;
      _tmp_918 <= 0;
      _tmp_919 <= 0;
      _tmp_920 <= 0;
      _tmp_921 <= 0;
      _tmp_922 <= 0;
      _tmp_923 <= 0;
      _tmp_924 <= 0;
      _tmp_925 <= 0;
      _tmp_926 <= 0;
      _tmp_927 <= 0;
      _tmp_928 <= 0;
      _tmp_929 <= 0;
      _tmp_930 <= 0;
      _tmp_931 <= 0;
      _tmp_932 <= 0;
      _tmp_933 <= 0;
      _tmp_934 <= 0;
      _mul_26_busy_reg <= 0;
    end else begin
      if(_mul_26_stream_oready) begin
        _mul_26_x_source_ram_renable <= 0;
        _mul_26_x_source_fifo_deq <= 0;
      end 
      _mul_26_x_idle <= _mul_26_x_idle;
      if(_mul_26_stream_oready) begin
        _mul_26_y_source_ram_renable <= 0;
        _mul_26_y_source_fifo_deq <= 0;
      end 
      _mul_26_y_idle <= _mul_26_y_idle;
      if(_mul_26_stream_oready) begin
        _mul_26_rshift_source_ram_renable <= 0;
        _mul_26_rshift_source_fifo_deq <= 0;
      end 
      _mul_26_rshift_idle <= _mul_26_rshift_idle;
      if(_mul_26_stream_oready) begin
        _mul_26_z_sink_wenable <= 0;
        _mul_26_z_sink_fifo_enq <= 0;
      end 
      if(_mul_26_stream_oready) begin
        __mul_26_stream_ivalid_1 <= _mul_26_stream_ivalid;
      end 
      if(_mul_26_stream_oready) begin
        __mul_26_stream_ivalid_2 <= __mul_26_stream_ivalid_1;
      end 
      if(_mul_26_stream_oready) begin
        __mul_26_stream_ivalid_3 <= __mul_26_stream_ivalid_2;
      end 
      if(_mul_26_stream_oready) begin
        __mul_26_stream_ivalid_4 <= __mul_26_stream_ivalid_3;
      end 
      if(_mul_26_stream_oready) begin
        __mul_26_stream_ivalid_5 <= __mul_26_stream_ivalid_4;
      end 
      if(_mul_26_stream_oready) begin
        __mul_26_stream_ivalid_6 <= __mul_26_stream_ivalid_5;
      end 
      if(_mul_26_stream_oready) begin
        __mul_26_stream_ivalid_7 <= __mul_26_stream_ivalid_6;
      end 
      if(_mul_26_stream_oready) begin
        __mul_26_stream_ivalid_8 <= __mul_26_stream_ivalid_7;
      end 
      if(_mul_26_stream_oready) begin
        _greaterthan_data_1523 <= mul_26_rshift_data > 1'sd0;
      end 
      if(_mul_26_stream_oready) begin
        _minus_data_1525 <= mul_26_rshift_data - 2'sd1;
      end 
      if(_mul_26_stream_oready) begin
        _greatereq_data_1536 <= mul_26_x_data >= 1'sd0;
      end 
      if(_mul_26_stream_oready) begin
        __delay_data_2082__variable_1520 <= mul_26_x_data;
      end 
      if(_mul_26_stream_oready) begin
        __delay_data_2085__variable_1521 <= mul_26_y_data;
      end 
      if(_mul_26_stream_oready) begin
        __delay_data_2088__variable_1522 <= mul_26_rshift_data;
      end 
      if(_mul_26_stream_oready) begin
        _sll_data_1527 <= 2'sd1 << _minus_data_1525;
      end 
      if(_mul_26_stream_oready) begin
        __delay_data_2079_greaterthan_1523 <= _greaterthan_data_1523;
      end 
      if(_mul_26_stream_oready) begin
        __delay_data_2080_greatereq_1536 <= _greatereq_data_1536;
      end 
      if(_mul_26_stream_oready) begin
        __delay_data_2083__delay_2082__variable_1520 <= __delay_data_2082__variable_1520;
      end 
      if(_mul_26_stream_oready) begin
        __delay_data_2086__delay_2085__variable_1521 <= __delay_data_2085__variable_1521;
      end 
      if(_mul_26_stream_oready) begin
        __delay_data_2089__delay_2088__variable_1522 <= __delay_data_2088__variable_1522;
      end 
      if(_mul_26_stream_oready) begin
        _cond_data_1533 <= (__delay_data_2079_greaterthan_1523)? _sll_data_1527 : 1'sd0;
      end 
      if(_mul_26_stream_oready) begin
        __delay_data_2081__delay_2080_greatereq_1536 <= __delay_data_2080_greatereq_1536;
      end 
      if(_mul_26_stream_oready) begin
        __delay_data_2084__delay_2083__delay_2082__variable_1520 <= __delay_data_2083__delay_2082__variable_1520;
      end 
      if(_mul_26_stream_oready) begin
        __delay_data_2087__delay_2086__delay_2085__variable_1521 <= __delay_data_2086__delay_2085__variable_1521;
      end 
      if(_mul_26_stream_oready) begin
        __delay_data_2090__delay_2089__delay_2088__variable_1522 <= __delay_data_2089__delay_2088__variable_1522;
      end 
      if(_mul_26_stream_oready) begin
        __muladd_madd_odata_reg_1539 <= __muladd_madd_odata_1539;
      end 
      if(_mul_26_stream_oready) begin
        __delay_data_2091__delay_2090__delay_2089____variable_1522 <= __delay_data_2090__delay_2089__delay_2088__variable_1522;
      end 
      if(_mul_26_stream_oready) begin
        __delay_data_2092__delay_2091__delay_2090____variable_1522 <= __delay_data_2091__delay_2090__delay_2089____variable_1522;
      end 
      if(_mul_26_stream_oready) begin
        __delay_data_2093__delay_2092__delay_2091____variable_1522 <= __delay_data_2092__delay_2091__delay_2090____variable_1522;
      end 
      if(_mul_26_stream_oready) begin
        __delay_data_2094__delay_2093__delay_2092____variable_1522 <= __delay_data_2093__delay_2092__delay_2091____variable_1522;
      end 
      if(_mul_26_stream_oready) begin
        _sra_data_1540 <= __muladd_data_1539 >>> __delay_data_2094__delay_2093__delay_2092____variable_1522;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_1520 <= _cond_data_1925;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_1521 <= __delay_data_2284_reinterpretcast_1889;
      end 
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        __variable_wdata_1522 <= _plus_data_2095;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_901 <= _mul_26_source_start;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_902 <= _tmp_901;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_903 <= _tmp_902;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_904 <= _mul_26_source_start;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_905 <= _tmp_904;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_906 <= _tmp_905;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_907 <= _tmp_906;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_908 <= _tmp_907;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_909 <= _tmp_908;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_910 <= _tmp_909;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_911 <= _tmp_910;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_912 <= _tmp_911;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_913 <= _tmp_912;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_914 <= _mul_26_source_stop;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_915 <= _tmp_914;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_916 <= _tmp_915;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_917 <= _tmp_916;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_918 <= _tmp_917;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_919 <= _tmp_918;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_920 <= _tmp_919;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_921 <= _tmp_920;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_922 <= _tmp_921;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_923 <= _tmp_922;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_924 <= _mul_26_source_busy;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_925 <= _tmp_924;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_926 <= _tmp_925;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_927 <= _tmp_926;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_928 <= _tmp_927;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_929 <= _tmp_928;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_930 <= _tmp_929;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_931 <= _tmp_930;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_932 <= _tmp_931;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_933 <= _tmp_932;
      end 
      if(_mul_26_stream_oready) begin
        _tmp_934 <= _mul_26_sink_busy;
      end 
      if(!_mul_26_sink_busy && _tmp_934) begin
        _mul_26_busy_reg <= 0;
      end 
      if(_mul_26_source_busy) begin
        _mul_26_busy_reg <= 1;
      end 
    end
  end

  localparam _mul_26_fsm_1 = 1;
  localparam _mul_26_fsm_2 = 2;
  localparam _mul_26_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mul_26_fsm <= _mul_26_fsm_init;
      _mul_26_source_start <= 0;
      _mul_26_source_busy <= 0;
      _mul_26_stream_ivalid <= 0;
    end else begin
      if(__stream_conv2d_4_stream_ivalid_1 && _stream_conv2d_4_stream_oready) begin
        _mul_26_stream_ivalid <= 1'd1;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_busy) begin
        _mul_26_source_busy <= _stream_conv2d_4_source_busy;
      end 
      if(_mul_26_stream_oready && _tmp_903) begin
        _mul_26_stream_ivalid <= 1;
      end 
      if(_mul_26_stream_oready && 1'd0) begin
        _mul_26_stream_ivalid <= 0;
      end 
      case(_mul_26_fsm)
        _mul_26_fsm_init: begin
          if(_mul_26_run_flag) begin
            _mul_26_source_start <= 1;
          end 
          if(_mul_26_run_flag) begin
            _mul_26_fsm <= _mul_26_fsm_1;
          end 
        end
        _mul_26_fsm_1: begin
          if(_mul_26_source_start && _mul_26_stream_oready) begin
            _mul_26_source_start <= 0;
            _mul_26_source_busy <= 1;
          end 
          if(_mul_26_source_start && _mul_26_stream_oready) begin
            _mul_26_fsm <= _mul_26_fsm_2;
          end 
        end
        _mul_26_fsm_2: begin
          if(_mul_26_stream_oready) begin
            _mul_26_fsm <= _mul_26_fsm_3;
          end 
        end
        _mul_26_fsm_3: begin
          if(_mul_26_stream_oready && 1'd0) begin
            _mul_26_source_busy <= 0;
          end 
          if(_mul_26_stream_oready && 1'd0 && _mul_26_run_flag) begin
            _mul_26_source_start <= 1;
          end 
          if(_mul_26_stream_oready && 1'd0) begin
            _mul_26_fsm <= _mul_26_fsm_init;
          end 
          if(_mul_26_stream_oready && 1'd0 && _mul_26_run_flag) begin
            _mul_26_fsm <= _mul_26_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __reduce_max_27_x_source_ram_renable <= 0;
      __reduce_max_27_x_source_fifo_deq <= 0;
      __reduce_max_27_x_idle <= 1;
      __reduce_max_27_data_sink_wenable <= 0;
      __reduce_max_27_data_sink_fifo_enq <= 0;
      __reduce_max_27_valid_sink_wenable <= 0;
      __reduce_max_27_valid_sink_fifo_enq <= 0;
      ___reduce_max_27_stream_ivalid_1 <= 0;
      _reducemax_data_1544 <= -17'sd32768;
      _reducemax_count_1544 <= 0;
      _reducemax_prev_count_max_1544 <= 0;
      _pulse_data_1546 <= 1'sd0;
      _pulse_count_1546 <= 0;
      _pulse_prev_count_max_1546 <= 0;
      __variable_wdata_1543 <= 0;
      __variable_wdata_1541 <= 0;
      __variable_wdata_1542 <= 0;
      _tmp_1235 <= 0;
      _tmp_1236 <= 0;
      _tmp_1237 <= 0;
      _tmp_1238 <= 0;
      _tmp_1239 <= 0;
      _tmp_1240 <= 0;
      _tmp_1241 <= 0;
      _tmp_1242 <= 0;
      _tmp_1243 <= 0;
      _tmp_1244 <= 0;
      _tmp_1245 <= 0;
      _tmp_1246 <= 0;
      _tmp_1247 <= 0;
      _tmp_1248 <= 0;
      _tmp_1249 <= 0;
      _tmp_1250 <= 0;
      _tmp_1251 <= 0;
      _tmp_1252 <= 0;
      _tmp_1253 <= 0;
      _tmp_1254 <= 0;
      __reduce_max_27_busy_reg <= 0;
    end else begin
      if(__reduce_max_27_stream_oready) begin
        __reduce_max_27_x_source_ram_renable <= 0;
        __reduce_max_27_x_source_fifo_deq <= 0;
      end 
      __reduce_max_27_x_idle <= __reduce_max_27_x_idle;
      if(__reduce_max_27_stream_oready) begin
        __reduce_max_27_data_sink_wenable <= 0;
        __reduce_max_27_data_sink_fifo_enq <= 0;
      end 
      if(__reduce_max_27_stream_oready) begin
        __reduce_max_27_valid_sink_wenable <= 0;
        __reduce_max_27_valid_sink_fifo_enq <= 0;
      end 
      if(__reduce_max_27_stream_oready) begin
        ___reduce_max_27_stream_ivalid_1 <= __reduce_max_27_stream_ivalid;
      end 
      if(__reduce_max_27_stream_ivalid && __reduce_max_27_stream_oready && _reducemax_reset_cond_1544) begin
        _reducemax_data_1544 <= -17'sd32768;
      end 
      if(__reduce_max_27_stream_ivalid && __reduce_max_27_stream_oready) begin
        _reducemax_count_1544 <= (_reducemax_current_count_1544 >= _reduce_max_27_size_data - 1)? 0 : _reducemax_current_count_1544 + 1;
      end 
      if(__reduce_max_27_stream_ivalid && __reduce_max_27_stream_oready) begin
        _reducemax_prev_count_max_1544 <= _reducemax_current_count_1544 >= _reduce_max_27_size_data - 1;
      end 
      if(__reduce_max_27_stream_ivalid && __reduce_max_27_stream_oready) begin
        _reducemax_data_1544 <= (_reducemax_current_data_1544 < _reduce_max_27_x_data)? _reduce_max_27_x_data : _reducemax_current_data_1544;
      end 
      if(__reduce_max_27_stream_ivalid && __reduce_max_27_stream_oready && _pulse_reset_cond_1546) begin
        _pulse_data_1546 <= 1'sd0;
      end 
      if(__reduce_max_27_stream_ivalid && __reduce_max_27_stream_oready) begin
        _pulse_count_1546 <= (_pulse_current_count_1546 >= _reduce_max_27_size_data - 1)? 0 : _pulse_current_count_1546 + 1;
      end 
      if(__reduce_max_27_stream_ivalid && __reduce_max_27_stream_oready) begin
        _pulse_prev_count_max_1546 <= _pulse_current_count_1546 >= _reduce_max_27_size_data - 1;
      end 
      if(__reduce_max_27_stream_ivalid && __reduce_max_27_stream_oready) begin
        _pulse_data_1546 <= _pulse_current_count_1546 >= _reduce_max_27_size_data - 1;
      end 
      if(__stream_max_pool_serial_6_stream_ivalid_3 && _stream_max_pool_serial_6_stream_oready) begin
        __variable_wdata_1543 <= __delay_data_2399__delay_2398__delay_2397__variable_2140;
      end 
      if(__stream_max_pool_serial_6_stream_ivalid_3 && _stream_max_pool_serial_6_stream_oready) begin
        __variable_wdata_1541 <= _cond_data_2151;
      end 
      if(__stream_max_pool_serial_6_stream_ivalid_3 && _stream_max_pool_serial_6_stream_oready) begin
        __variable_wdata_1542 <= __delay_data_2402__delay_2401__delay_2400__variable_2137;
      end 
      if(__reduce_max_27_stream_oready) begin
        _tmp_1235 <= __reduce_max_27_source_start;
      end 
      if(__reduce_max_27_stream_oready) begin
        _tmp_1236 <= _tmp_1235;
      end 
      if(__reduce_max_27_stream_oready) begin
        _tmp_1237 <= _tmp_1236;
      end 
      if(__reduce_max_27_stream_oready) begin
        _tmp_1238 <= __reduce_max_27_source_start;
      end 
      if(__reduce_max_27_stream_oready) begin
        _tmp_1239 <= _tmp_1238;
      end 
      if(__reduce_max_27_stream_oready) begin
        _tmp_1240 <= _tmp_1239;
      end 
      if(__reduce_max_27_stream_oready && _tmp_1240) begin
        __variable_wdata_1543 <= 1;
      end 
      if(__reduce_max_27_stream_oready) begin
        _tmp_1241 <= __reduce_max_27_source_start;
      end 
      if(__reduce_max_27_stream_oready) begin
        _tmp_1242 <= _tmp_1241;
      end 
      if(__reduce_max_27_stream_oready) begin
        _tmp_1243 <= _tmp_1242;
      end 
      if(__reduce_max_27_stream_oready) begin
        _tmp_1244 <= _tmp_1243;
      end 
      if(__reduce_max_27_stream_oready && _tmp_1244) begin
        __variable_wdata_1543 <= 0;
      end 
      if(__reduce_max_27_stream_oready && 1'd0) begin
        __variable_wdata_1543 <= 1;
      end 
      if(__reduce_max_27_stream_oready) begin
        _tmp_1245 <= __reduce_max_27_source_start;
      end 
      if(__reduce_max_27_stream_oready) begin
        _tmp_1246 <= _tmp_1245;
      end 
      if(__reduce_max_27_stream_oready) begin
        _tmp_1247 <= _tmp_1246;
      end 
      if(__reduce_max_27_stream_oready) begin
        _tmp_1248 <= __reduce_max_27_source_stop;
      end 
      if(__reduce_max_27_stream_oready) begin
        _tmp_1249 <= _tmp_1248;
      end 
      if(__reduce_max_27_stream_oready) begin
        _tmp_1250 <= _tmp_1249;
      end 
      if(__reduce_max_27_stream_oready) begin
        _tmp_1251 <= __reduce_max_27_source_busy;
      end 
      if(__reduce_max_27_stream_oready) begin
        _tmp_1252 <= _tmp_1251;
      end 
      if(__reduce_max_27_stream_oready) begin
        _tmp_1253 <= _tmp_1252;
      end 
      if(__reduce_max_27_stream_oready) begin
        _tmp_1254 <= __reduce_max_27_sink_busy;
      end 
      if(!__reduce_max_27_sink_busy && _tmp_1254) begin
        __reduce_max_27_busy_reg <= 0;
      end 
      if(__reduce_max_27_source_busy) begin
        __reduce_max_27_busy_reg <= 1;
      end 
    end
  end

  localparam __reduce_max_27_fsm_1 = 1;
  localparam __reduce_max_27_fsm_2 = 2;
  localparam __reduce_max_27_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      __reduce_max_27_fsm <= __reduce_max_27_fsm_init;
      __reduce_max_27_source_start <= 0;
      __reduce_max_27_source_busy <= 0;
      __reduce_max_27_stream_ivalid <= 0;
    end else begin
      if(__stream_max_pool_serial_6_stream_ivalid_3 && _stream_max_pool_serial_6_stream_oready) begin
        __reduce_max_27_stream_ivalid <= 1'd1;
      end 
      if(_stream_max_pool_serial_6_stream_oready && _stream_max_pool_serial_6_busy) begin
        __reduce_max_27_source_busy <= _stream_max_pool_serial_6_source_busy;
      end 
      if(__reduce_max_27_stream_oready && _tmp_1237) begin
        __reduce_max_27_stream_ivalid <= 1;
      end 
      if(__reduce_max_27_stream_oready && 1'd0) begin
        __reduce_max_27_stream_ivalid <= 0;
      end 
      case(__reduce_max_27_fsm)
        __reduce_max_27_fsm_init: begin
          if(__reduce_max_27_run_flag) begin
            __reduce_max_27_source_start <= 1;
          end 
          if(__reduce_max_27_run_flag) begin
            __reduce_max_27_fsm <= __reduce_max_27_fsm_1;
          end 
        end
        __reduce_max_27_fsm_1: begin
          if(__reduce_max_27_source_start && __reduce_max_27_stream_oready) begin
            __reduce_max_27_source_start <= 0;
            __reduce_max_27_source_busy <= 1;
          end 
          if(__reduce_max_27_source_start && __reduce_max_27_stream_oready) begin
            __reduce_max_27_fsm <= __reduce_max_27_fsm_2;
          end 
        end
        __reduce_max_27_fsm_2: begin
          if(__reduce_max_27_stream_oready) begin
            __reduce_max_27_fsm <= __reduce_max_27_fsm_3;
          end 
        end
        __reduce_max_27_fsm_3: begin
          if(__reduce_max_27_stream_oready && 1'd0) begin
            __reduce_max_27_source_busy <= 0;
          end 
          if(__reduce_max_27_stream_oready && 1'd0 && __reduce_max_27_run_flag) begin
            __reduce_max_27_source_start <= 1;
          end 
          if(__reduce_max_27_stream_oready && 1'd0) begin
            __reduce_max_27_fsm <= __reduce_max_27_fsm_init;
          end 
          if(__reduce_max_27_stream_oready && 1'd0 && __reduce_max_27_run_flag) begin
            __reduce_max_27_fsm <= __reduce_max_27_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_7_source_ram_renable <= 0;
      _stream_conv2d_4_source_7_source_fifo_deq <= 0;
      _stream_conv2d_4_source_7_idle <= 1;
      _stream_conv2d_4_source_9_source_ram_renable <= 0;
      _stream_conv2d_4_source_9_source_fifo_deq <= 0;
      _stream_conv2d_4_source_9_idle <= 1;
      _stream_conv2d_4_source_11_source_ram_renable <= 0;
      _stream_conv2d_4_source_11_source_fifo_deq <= 0;
      _stream_conv2d_4_source_11_idle <= 1;
      _stream_conv2d_4_source_13_source_ram_renable <= 0;
      _stream_conv2d_4_source_13_source_fifo_deq <= 0;
      _stream_conv2d_4_source_13_idle <= 1;
      _stream_conv2d_4_source_15_source_ram_renable <= 0;
      _stream_conv2d_4_source_15_source_fifo_deq <= 0;
      _stream_conv2d_4_source_15_idle <= 1;
      _stream_conv2d_4_source_20_source_ram_renable <= 0;
      _stream_conv2d_4_source_20_source_fifo_deq <= 0;
      _stream_conv2d_4_source_20_idle <= 1;
      _stream_conv2d_4_source_21_source_ram_renable <= 0;
      _stream_conv2d_4_source_21_source_fifo_deq <= 0;
      _stream_conv2d_4_source_21_idle <= 1;
      _stream_conv2d_4_source_22_source_ram_renable <= 0;
      _stream_conv2d_4_source_22_source_fifo_deq <= 0;
      _stream_conv2d_4_source_22_idle <= 1;
      _stream_conv2d_4_source_23_source_ram_renable <= 0;
      _stream_conv2d_4_source_23_source_fifo_deq <= 0;
      _stream_conv2d_4_source_23_idle <= 1;
      _stream_conv2d_4_source_24_source_ram_renable <= 0;
      _stream_conv2d_4_source_24_source_fifo_deq <= 0;
      _stream_conv2d_4_source_24_idle <= 1;
      _stream_conv2d_4_source_25_source_ram_renable <= 0;
      _stream_conv2d_4_source_25_source_fifo_deq <= 0;
      _stream_conv2d_4_source_25_idle <= 1;
      _stream_conv2d_4_source_26_source_ram_renable <= 0;
      _stream_conv2d_4_source_26_source_fifo_deq <= 0;
      _stream_conv2d_4_source_26_idle <= 1;
      _stream_conv2d_4_source_27_source_ram_renable <= 0;
      _stream_conv2d_4_source_27_source_fifo_deq <= 0;
      _stream_conv2d_4_source_27_idle <= 1;
      _stream_conv2d_4_source_28_source_ram_renable <= 0;
      _stream_conv2d_4_source_28_source_fifo_deq <= 0;
      _stream_conv2d_4_source_28_idle <= 1;
      _stream_conv2d_4_source_29_source_ram_renable <= 0;
      _stream_conv2d_4_source_29_source_fifo_deq <= 0;
      _stream_conv2d_4_source_29_idle <= 1;
      _stream_conv2d_4_source_30_source_ram_renable <= 0;
      _stream_conv2d_4_source_30_source_fifo_deq <= 0;
      _stream_conv2d_4_source_30_idle <= 1;
      _stream_conv2d_4_source_31_source_ram_renable <= 0;
      _stream_conv2d_4_source_31_source_fifo_deq <= 0;
      _stream_conv2d_4_source_31_idle <= 1;
      _stream_conv2d_4_source_32_source_ram_renable <= 0;
      _stream_conv2d_4_source_32_source_fifo_deq <= 0;
      _stream_conv2d_4_source_32_idle <= 1;
      _stream_conv2d_4_source_33_source_ram_renable <= 0;
      _stream_conv2d_4_source_33_source_fifo_deq <= 0;
      _stream_conv2d_4_source_33_idle <= 1;
      _stream_conv2d_4_source_34_source_ram_renable <= 0;
      _stream_conv2d_4_source_34_source_fifo_deq <= 0;
      _stream_conv2d_4_source_34_idle <= 1;
      _stream_conv2d_4_source_35_source_ram_renable <= 0;
      _stream_conv2d_4_source_35_source_fifo_deq <= 0;
      _stream_conv2d_4_source_35_idle <= 1;
      _stream_conv2d_4_source_36_source_ram_renable <= 0;
      _stream_conv2d_4_source_36_source_fifo_deq <= 0;
      _stream_conv2d_4_source_36_idle <= 1;
      _stream_conv2d_4_source_37_source_ram_renable <= 0;
      _stream_conv2d_4_source_37_source_fifo_deq <= 0;
      _stream_conv2d_4_source_37_idle <= 1;
      _stream_conv2d_4_sink_50_sink_wenable <= 0;
      _stream_conv2d_4_sink_50_sink_fifo_enq <= 0;
      _stream_conv2d_4_sink_51_sink_wenable <= 0;
      _stream_conv2d_4_sink_51_sink_fifo_enq <= 0;
      __stream_conv2d_4_stream_ivalid_1 <= 0;
      __stream_conv2d_4_stream_ivalid_2 <= 0;
      __stream_conv2d_4_stream_ivalid_3 <= 0;
      __stream_conv2d_4_stream_ivalid_4 <= 0;
      __stream_conv2d_4_stream_ivalid_5 <= 0;
      __stream_conv2d_4_stream_ivalid_6 <= 0;
      __stream_conv2d_4_stream_ivalid_7 <= 0;
      __stream_conv2d_4_stream_ivalid_8 <= 0;
      __stream_conv2d_4_stream_ivalid_9 <= 0;
      __stream_conv2d_4_stream_ivalid_10 <= 0;
      __stream_conv2d_4_stream_ivalid_11 <= 0;
      __stream_conv2d_4_stream_ivalid_12 <= 0;
      __stream_conv2d_4_stream_ivalid_13 <= 0;
      __stream_conv2d_4_stream_ivalid_14 <= 0;
      __stream_conv2d_4_stream_ivalid_15 <= 0;
      __stream_conv2d_4_stream_ivalid_16 <= 0;
      __stream_conv2d_4_stream_ivalid_17 <= 0;
      __stream_conv2d_4_stream_ivalid_18 <= 0;
      __stream_conv2d_4_stream_ivalid_19 <= 0;
      __stream_conv2d_4_stream_ivalid_20 <= 0;
      __stream_conv2d_4_stream_ivalid_21 <= 0;
      __stream_conv2d_4_stream_ivalid_22 <= 0;
      __stream_conv2d_4_stream_ivalid_23 <= 0;
      __stream_conv2d_4_stream_ivalid_24 <= 0;
      __stream_conv2d_4_stream_ivalid_25 <= 0;
      __stream_conv2d_4_stream_ivalid_26 <= 0;
      __stream_conv2d_4_stream_ivalid_27 <= 0;
      __stream_conv2d_4_stream_ivalid_28 <= 0;
      __stream_conv2d_4_stream_ivalid_29 <= 0;
      __stream_conv2d_4_stream_ivalid_30 <= 0;
      __stream_conv2d_4_stream_ivalid_31 <= 0;
      _eq_data_1611 <= 0;
      _eq_data_1615 <= 0;
      _eq_data_1618 <= 0;
      _eq_data_1621 <= 0;
      _eq_data_1625 <= 0;
      _eq_data_1628 <= 0;
      _eq_data_1631 <= 0;
      _eq_data_1635 <= 0;
      _eq_data_1638 <= 0;
      _eq_data_1641 <= 0;
      _eq_data_1645 <= 0;
      _eq_data_1648 <= 0;
      _eq_data_1651 <= 0;
      _eq_data_1655 <= 0;
      _eq_data_1658 <= 0;
      _eq_data_1661 <= 0;
      _eq_data_1665 <= 0;
      _eq_data_1668 <= 0;
      _eq_data_1671 <= 0;
      _eq_data_1675 <= 0;
      _eq_data_1678 <= 0;
      _eq_data_1681 <= 0;
      _eq_data_1685 <= 0;
      _eq_data_1688 <= 0;
      _eq_data_1691 <= 0;
      _eq_data_1695 <= 0;
      _eq_data_1698 <= 0;
      _eq_data_1701 <= 0;
      _eq_data_1705 <= 0;
      _eq_data_1708 <= 0;
      _eq_data_1711 <= 0;
      _eq_data_1715 <= 0;
      _eq_data_1718 <= 0;
      _eq_data_1721 <= 0;
      _eq_data_1725 <= 0;
      _eq_data_1728 <= 0;
      _eq_data_1731 <= 0;
      _eq_data_1735 <= 0;
      _eq_data_1738 <= 0;
      _eq_data_1741 <= 0;
      _eq_data_1745 <= 0;
      _eq_data_1748 <= 0;
      _eq_data_1751 <= 0;
      _eq_data_1755 <= 0;
      _eq_data_1758 <= 0;
      _eq_data_1761 <= 0;
      _eq_data_1765 <= 0;
      _eq_data_1768 <= 0;
      _eq_data_1771 <= 0;
      _eq_data_1775 <= 0;
      _eq_data_1778 <= 0;
      _eq_data_1781 <= 0;
      _eq_data_1785 <= 0;
      _eq_data_1788 <= 0;
      _plus_data_1943 <= 0;
      _plus_data_1962 <= 0;
      _plus_data_1981 <= 0;
      _plus_data_2000 <= 0;
      _plus_data_2019 <= 0;
      _plus_data_2038 <= 0;
      _plus_data_2057 <= 0;
      _plus_data_2076 <= 0;
      _plus_data_2095 <= 0;
      _plus_data_2111 <= 0;
      _plus_data_2130 <= 0;
      __delay_data_2258__variable_1604 <= 0;
      __delay_data_2259__variable_1603 <= 0;
      __delay_data_2260__variable_1602 <= 0;
      __delay_data_2261__variable_1607 <= 0;
      __delay_data_2262__variable_1606 <= 0;
      __delay_data_2263__variable_1605 <= 0;
      __delay_data_2264__variable_1610 <= 0;
      __delay_data_2265__variable_1609 <= 0;
      __delay_data_2266__variable_1608 <= 0;
      __delay_data_2267_pointer_1890 <= 0;
      __delay_data_2268_reinterpretcast_1881 <= 0;
      __delay_data_2269_pointer_1892 <= 0;
      __delay_data_2270_reinterpretcast_1882 <= 0;
      __delay_data_2271_pointer_1894 <= 0;
      __delay_data_2272_reinterpretcast_1883 <= 0;
      __delay_data_2273_pointer_1896 <= 0;
      __delay_data_2274_reinterpretcast_1884 <= 0;
      __delay_data_2275_pointer_1898 <= 0;
      __delay_data_2276_reinterpretcast_1885 <= 0;
      __delay_data_2277_pointer_1900 <= 0;
      __delay_data_2278_reinterpretcast_1886 <= 0;
      __delay_data_2279_pointer_1902 <= 0;
      __delay_data_2280_reinterpretcast_1887 <= 0;
      __delay_data_2281_pointer_1904 <= 0;
      __delay_data_2282_reinterpretcast_1888 <= 0;
      __delay_data_2283_pointer_1906 <= 0;
      __delay_data_2284_reinterpretcast_1889 <= 0;
      __delay_data_2285__variable_1553 <= 0;
      __delay_data_2310__variable_1548 <= 0;
      __delay_data_2323_cond_1569 <= 0;
      __delay_data_2342_cond_1576 <= 0;
      __delay_data_2286__delay_2285__variable_1553 <= 0;
      __delay_data_2298_plus_2111 <= 0;
      __delay_data_2311__delay_2310__variable_1548 <= 0;
      __delay_data_2324__delay_2323_cond_1569 <= 0;
      __delay_data_2343__delay_2342_cond_1576 <= 0;
      __delay_data_2362_plus_2130 <= 0;
      __delay_data_2287__delay_2286__delay_2285__variable_1553 <= 0;
      __delay_data_2299__delay_2298_plus_2111 <= 0;
      __delay_data_2312__delay_2311__delay_2310__variable_1548 <= 0;
      __delay_data_2325__delay_2324__delay_2323_cond_1569 <= 0;
      __delay_data_2344__delay_2343__delay_2342_cond_1576 <= 0;
      __delay_data_2363__delay_2362_plus_2130 <= 0;
      __delay_data_2288__delay_2287__delay_2286____variable_1553 <= 0;
      __delay_data_2300__delay_2299__delay_2298_plus_2111 <= 0;
      __delay_data_2313__delay_2312__delay_2311____variable_1548 <= 0;
      __delay_data_2326__delay_2325__delay_2324___cond_1569 <= 0;
      __delay_data_2345__delay_2344__delay_2343___cond_1576 <= 0;
      __delay_data_2364__delay_2363__delay_2362_plus_2130 <= 0;
      __delay_data_2289__delay_2288__delay_2287____variable_1553 <= 0;
      __delay_data_2301__delay_2300__delay_2299___plus_2111 <= 0;
      __delay_data_2314__delay_2313__delay_2312____variable_1548 <= 0;
      __delay_data_2327__delay_2326__delay_2325___cond_1569 <= 0;
      __delay_data_2346__delay_2345__delay_2344___cond_1576 <= 0;
      __delay_data_2365__delay_2364__delay_2363___plus_2130 <= 0;
      __delay_data_2290__delay_2289__delay_2288____variable_1553 <= 0;
      __delay_data_2302__delay_2301__delay_2300___plus_2111 <= 0;
      __delay_data_2315__delay_2314__delay_2313____variable_1548 <= 0;
      __delay_data_2328__delay_2327__delay_2326___cond_1569 <= 0;
      __delay_data_2347__delay_2346__delay_2345___cond_1576 <= 0;
      __delay_data_2366__delay_2365__delay_2364___plus_2130 <= 0;
      __delay_data_2291__delay_2290__delay_2289____variable_1553 <= 0;
      __delay_data_2303__delay_2302__delay_2301___plus_2111 <= 0;
      __delay_data_2316__delay_2315__delay_2314____variable_1548 <= 0;
      __delay_data_2329__delay_2328__delay_2327___cond_1569 <= 0;
      __delay_data_2348__delay_2347__delay_2346___cond_1576 <= 0;
      __delay_data_2367__delay_2366__delay_2365___plus_2130 <= 0;
      __delay_data_2292__delay_2291__delay_2290____variable_1553 <= 0;
      __delay_data_2304__delay_2303__delay_2302___plus_2111 <= 0;
      __delay_data_2317__delay_2316__delay_2315____variable_1548 <= 0;
      __delay_data_2330__delay_2329__delay_2328___cond_1569 <= 0;
      __delay_data_2349__delay_2348__delay_2347___cond_1576 <= 0;
      __delay_data_2368__delay_2367__delay_2366___plus_2130 <= 0;
      __delay_data_2293__delay_2292__delay_2291____variable_1553 <= 0;
      __delay_data_2305__delay_2304__delay_2303___plus_2111 <= 0;
      __delay_data_2318__delay_2317__delay_2316____variable_1548 <= 0;
      __delay_data_2331__delay_2330__delay_2329___cond_1569 <= 0;
      __delay_data_2350__delay_2349__delay_2348___cond_1576 <= 0;
      __delay_data_2369__delay_2368__delay_2367___plus_2130 <= 0;
      __delay_data_2294__delay_2293__delay_2292____variable_1553 <= 0;
      __delay_data_2306__delay_2305__delay_2304___plus_2111 <= 0;
      __delay_data_2319__delay_2318__delay_2317____variable_1548 <= 0;
      __delay_data_2332__delay_2331__delay_2330___cond_1569 <= 0;
      __delay_data_2351__delay_2350__delay_2349___cond_1576 <= 0;
      __delay_data_2370__delay_2369__delay_2368___plus_2130 <= 0;
      __delay_data_2295__delay_2294__delay_2293____variable_1553 <= 0;
      __delay_data_2307__delay_2306__delay_2305___plus_2111 <= 0;
      __delay_data_2320__delay_2319__delay_2318____variable_1548 <= 0;
      __delay_data_2333__delay_2332__delay_2331___cond_1569 <= 0;
      __delay_data_2352__delay_2351__delay_2350___cond_1576 <= 0;
      __delay_data_2371__delay_2370__delay_2369___plus_2130 <= 0;
      __delay_data_2296__delay_2295__delay_2294____variable_1553 <= 0;
      __delay_data_2308__delay_2307__delay_2306___plus_2111 <= 0;
      __delay_data_2321__delay_2320__delay_2319____variable_1548 <= 0;
      __delay_data_2334__delay_2333__delay_2332___cond_1569 <= 0;
      __delay_data_2353__delay_2352__delay_2351___cond_1576 <= 0;
      __delay_data_2372__delay_2371__delay_2370___plus_2130 <= 0;
      __delay_data_2297__delay_2296__delay_2295____variable_1553 <= 0;
      __delay_data_2309__delay_2308__delay_2307___plus_2111 <= 0;
      __delay_data_2322__delay_2321__delay_2320____variable_1548 <= 0;
      __delay_data_2335__delay_2334__delay_2333___cond_1569 <= 0;
      __delay_data_2354__delay_2353__delay_2352___cond_1576 <= 0;
      __delay_data_2373__delay_2372__delay_2371___plus_2130 <= 0;
      __delay_data_2336__delay_2335__delay_2334___cond_1569 <= 0;
      __delay_data_2355__delay_2354__delay_2353___cond_1576 <= 0;
      __delay_data_2374__delay_2373__delay_2372___plus_2130 <= 0;
      __delay_data_2337__delay_2336__delay_2335___cond_1569 <= 0;
      __delay_data_2356__delay_2355__delay_2354___cond_1576 <= 0;
      __delay_data_2375__delay_2374__delay_2373___plus_2130 <= 0;
      __delay_data_2338__delay_2337__delay_2336___cond_1569 <= 0;
      __delay_data_2357__delay_2356__delay_2355___cond_1576 <= 0;
      __delay_data_2376__delay_2375__delay_2374___plus_2130 <= 0;
      __delay_data_2339__delay_2338__delay_2337___cond_1569 <= 0;
      __delay_data_2358__delay_2357__delay_2356___cond_1576 <= 0;
      __delay_data_2377__delay_2376__delay_2375___plus_2130 <= 0;
      __delay_data_2340__delay_2339__delay_2338___cond_1569 <= 0;
      __delay_data_2359__delay_2358__delay_2357___cond_1576 <= 0;
      __delay_data_2378__delay_2377__delay_2376___plus_2130 <= 0;
      __delay_data_2341__delay_2340__delay_2339___cond_1569 <= 0;
      __delay_data_2360__delay_2359__delay_2358___cond_1576 <= 0;
      __delay_data_2379__delay_2378__delay_2377___plus_2130 <= 0;
      _plus_data_2114 <= 0;
      __delay_data_2361__delay_2360__delay_2359___cond_1576 <= 0;
      __delay_data_2380__delay_2379__delay_2378___plus_2130 <= 0;
      __delay_data_2382__substreamoutput_2113 <= 0;
      __delay_data_2383__delay_2382__substreamoutput_2113 <= 0;
      __delay_data_2384__delay_2383____substreamoutput_2113 <= 0;
      __delay_data_2385__delay_2384____substreamoutput_2113 <= 0;
      __delay_data_2386__delay_2385____substreamoutput_2113 <= 0;
      __delay_data_2387__delay_2386____substreamoutput_2113 <= 0;
      __delay_data_2388__delay_2387____substreamoutput_2113 <= 0;
      __delay_data_2389__delay_2388____substreamoutput_2113 <= 0;
      __delay_data_2390__delay_2389____substreamoutput_2113 <= 0;
      __delay_data_2391__delay_2390____substreamoutput_2113 <= 0;
      _greaterthan_data_2133 <= 0;
      __delay_data_2381__substreamoutput_2131 <= 0;
      __delay_data_2392__delay_2391____substreamoutput_2113 <= 0;
      _cond_data_2135 <= 0;
      __delay_data_2393__delay_2392____substreamoutput_2113 <= 0;
      _stream_conv2d_4_parameter_0_next_parameter_data <= 0;
      __variable_wdata_1548 <= 0;
      _stream_conv2d_4_parameter_1_next_parameter_data <= 0;
      __variable_wdata_1549 <= 0;
      _stream_conv2d_4_parameter_2_next_parameter_data <= 0;
      __variable_wdata_1550 <= 0;
      _stream_conv2d_4_parameter_3_next_parameter_data <= 0;
      __variable_wdata_1551 <= 0;
      _stream_conv2d_4_parameter_4_next_parameter_data <= 0;
      __variable_wdata_1552 <= 0;
      _stream_conv2d_4_parameter_6_next_parameter_data <= 0;
      __variable_wdata_1563 <= 0;
      _stream_conv2d_4_source_7_source_mode <= 5'b0;
      _stream_conv2d_4_source_7_source_offset <= 0;
      _source_stream_conv2d_4_source_7_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_7_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_7_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_7_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_7_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_7_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_7_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_7_pat_stride_3 <= 0;
      _stream_conv2d_4_source_7_source_sel <= 0;
      _stream_conv2d_4_source_7_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_7_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_7_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_7_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_7_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_7_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_7_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_7_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_7_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_7_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_7_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_7_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_7_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_7_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_7_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_7_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_7_pat_stride_buf_3 <= 0;
      __variable_wdata_1564 <= 0;
      _stream_conv2d_4_source_7_source_ram_raddr <= 0;
      _stream_conv2d_4_parameter_8_next_parameter_data <= 0;
      __variable_wdata_1570 <= 0;
      _stream_conv2d_4_source_9_source_mode <= 5'b0;
      _stream_conv2d_4_source_9_source_offset <= 0;
      _source_stream_conv2d_4_source_9_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_9_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_9_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_9_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_9_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_9_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_9_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_9_pat_stride_3 <= 0;
      _stream_conv2d_4_source_9_source_sel <= 0;
      _stream_conv2d_4_source_9_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_9_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_9_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_9_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_9_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_9_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_9_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_9_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_9_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_9_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_9_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_9_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_9_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_9_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_9_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_9_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_9_pat_stride_buf_3 <= 0;
      __variable_wdata_1571 <= 0;
      _stream_conv2d_4_source_9_source_ram_raddr <= 0;
      _stream_conv2d_4_parameter_10_next_parameter_data <= 0;
      __variable_wdata_1577 <= 0;
      _stream_conv2d_4_source_11_source_mode <= 5'b0;
      _stream_conv2d_4_source_11_source_empty_data <= 0;
      __variable_wdata_1578 <= 0;
      _stream_conv2d_4_parameter_12_next_parameter_data <= 0;
      __variable_wdata_1584 <= 0;
      _stream_conv2d_4_source_13_source_mode <= 5'b0;
      _stream_conv2d_4_source_13_source_empty_data <= 0;
      __variable_wdata_1585 <= 0;
      _stream_conv2d_4_parameter_14_next_parameter_data <= 0;
      __variable_wdata_1591 <= 0;
      _stream_conv2d_4_source_15_source_mode <= 5'b0;
      _stream_conv2d_4_source_15_source_empty_data <= 0;
      __variable_wdata_1592 <= 0;
      _stream_conv2d_4_parameter_16_next_parameter_data <= 0;
      __variable_wdata_1598 <= 0;
      _stream_conv2d_4_parameter_17_next_parameter_data <= 0;
      __variable_wdata_1599 <= 0;
      _stream_conv2d_4_parameter_18_next_parameter_data <= 0;
      __variable_wdata_1600 <= 0;
      _stream_conv2d_4_parameter_19_next_parameter_data <= 0;
      __variable_wdata_1601 <= 0;
      _stream_conv2d_4_source_20_source_mode <= 5'b0;
      _stream_conv2d_4_source_20_source_offset <= 0;
      _source_stream_conv2d_4_source_20_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_20_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_20_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_20_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_20_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_20_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_20_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_20_pat_stride_3 <= 0;
      _stream_conv2d_4_source_20_source_sel <= 0;
      _stream_conv2d_4_source_20_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_20_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_20_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_20_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_20_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_20_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_20_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_20_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_20_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_20_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_20_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_20_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_20_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_20_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_20_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_20_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_20_pat_stride_buf_3 <= 0;
      __variable_wdata_1602 <= 0;
      _stream_conv2d_4_source_20_source_ram_raddr <= 0;
      _stream_conv2d_4_source_21_source_mode <= 5'b0;
      _stream_conv2d_4_source_21_source_offset <= 0;
      _source_stream_conv2d_4_source_21_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_21_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_21_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_21_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_21_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_21_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_21_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_21_pat_stride_3 <= 0;
      _stream_conv2d_4_source_21_source_sel <= 0;
      _stream_conv2d_4_source_21_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_21_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_21_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_21_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_21_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_21_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_21_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_21_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_21_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_21_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_21_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_21_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_21_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_21_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_21_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_21_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_21_pat_stride_buf_3 <= 0;
      __variable_wdata_1603 <= 0;
      _stream_conv2d_4_source_21_source_ram_raddr <= 0;
      _stream_conv2d_4_source_22_source_mode <= 5'b0;
      _stream_conv2d_4_source_22_source_offset <= 0;
      _source_stream_conv2d_4_source_22_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_22_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_22_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_22_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_22_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_22_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_22_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_22_pat_stride_3 <= 0;
      _stream_conv2d_4_source_22_source_sel <= 0;
      _stream_conv2d_4_source_22_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_22_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_22_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_22_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_22_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_22_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_22_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_22_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_22_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_22_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_22_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_22_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_22_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_22_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_22_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_22_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_22_pat_stride_buf_3 <= 0;
      __variable_wdata_1604 <= 0;
      _stream_conv2d_4_source_22_source_ram_raddr <= 0;
      _stream_conv2d_4_source_23_source_mode <= 5'b0;
      _stream_conv2d_4_source_23_source_offset <= 0;
      _source_stream_conv2d_4_source_23_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_23_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_23_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_23_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_23_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_23_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_23_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_23_pat_stride_3 <= 0;
      _stream_conv2d_4_source_23_source_sel <= 0;
      _stream_conv2d_4_source_23_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_23_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_23_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_23_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_23_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_23_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_23_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_23_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_23_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_23_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_23_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_23_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_23_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_23_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_23_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_23_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_23_pat_stride_buf_3 <= 0;
      __variable_wdata_1605 <= 0;
      _stream_conv2d_4_source_23_source_ram_raddr <= 0;
      _stream_conv2d_4_source_24_source_mode <= 5'b0;
      _stream_conv2d_4_source_24_source_offset <= 0;
      _source_stream_conv2d_4_source_24_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_24_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_24_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_24_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_24_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_24_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_24_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_24_pat_stride_3 <= 0;
      _stream_conv2d_4_source_24_source_sel <= 0;
      _stream_conv2d_4_source_24_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_24_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_24_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_24_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_24_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_24_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_24_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_24_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_24_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_24_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_24_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_24_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_24_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_24_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_24_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_24_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_24_pat_stride_buf_3 <= 0;
      __variable_wdata_1606 <= 0;
      _stream_conv2d_4_source_24_source_ram_raddr <= 0;
      _stream_conv2d_4_source_25_source_mode <= 5'b0;
      _stream_conv2d_4_source_25_source_offset <= 0;
      _source_stream_conv2d_4_source_25_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_25_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_25_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_25_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_25_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_25_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_25_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_25_pat_stride_3 <= 0;
      _stream_conv2d_4_source_25_source_sel <= 0;
      _stream_conv2d_4_source_25_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_25_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_25_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_25_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_25_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_25_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_25_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_25_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_25_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_25_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_25_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_25_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_25_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_25_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_25_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_25_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_25_pat_stride_buf_3 <= 0;
      __variable_wdata_1607 <= 0;
      _stream_conv2d_4_source_25_source_ram_raddr <= 0;
      _stream_conv2d_4_source_26_source_mode <= 5'b0;
      _stream_conv2d_4_source_26_source_offset <= 0;
      _source_stream_conv2d_4_source_26_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_26_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_26_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_26_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_26_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_26_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_26_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_26_pat_stride_3 <= 0;
      _stream_conv2d_4_source_26_source_sel <= 0;
      _stream_conv2d_4_source_26_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_26_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_26_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_26_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_26_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_26_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_26_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_26_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_26_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_26_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_26_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_26_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_26_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_26_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_26_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_26_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_26_pat_stride_buf_3 <= 0;
      __variable_wdata_1608 <= 0;
      _stream_conv2d_4_source_26_source_ram_raddr <= 0;
      _stream_conv2d_4_source_27_source_mode <= 5'b0;
      _stream_conv2d_4_source_27_source_offset <= 0;
      _source_stream_conv2d_4_source_27_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_27_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_27_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_27_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_27_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_27_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_27_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_27_pat_stride_3 <= 0;
      _stream_conv2d_4_source_27_source_sel <= 0;
      _stream_conv2d_4_source_27_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_27_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_27_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_27_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_27_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_27_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_27_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_27_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_27_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_27_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_27_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_27_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_27_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_27_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_27_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_27_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_27_pat_stride_buf_3 <= 0;
      __variable_wdata_1609 <= 0;
      _stream_conv2d_4_source_27_source_ram_raddr <= 0;
      _stream_conv2d_4_source_28_source_mode <= 5'b0;
      _stream_conv2d_4_source_28_source_offset <= 0;
      _source_stream_conv2d_4_source_28_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_28_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_28_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_28_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_28_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_28_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_28_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_28_pat_stride_3 <= 0;
      _stream_conv2d_4_source_28_source_sel <= 0;
      _stream_conv2d_4_source_28_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_28_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_28_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_28_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_28_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_28_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_28_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_28_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_28_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_28_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_28_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_28_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_28_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_28_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_28_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_28_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_28_pat_stride_buf_3 <= 0;
      __variable_wdata_1610 <= 0;
      _stream_conv2d_4_source_28_source_ram_raddr <= 0;
      _stream_conv2d_4_source_29_source_mode <= 5'b0;
      _stream_conv2d_4_source_29_source_offset <= 0;
      _source_stream_conv2d_4_source_29_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_29_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_29_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_29_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_29_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_29_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_29_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_29_pat_stride_3 <= 0;
      _stream_conv2d_4_source_29_source_sel <= 0;
      _stream_conv2d_4_source_29_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_29_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_29_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_29_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_29_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_29_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_29_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_29_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_29_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_29_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_29_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_29_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_29_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_29_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_29_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_29_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_29_pat_stride_buf_3 <= 0;
      __variable_wdata_1836 <= 0;
      _stream_conv2d_4_source_29_source_ram_raddr <= 0;
      _stream_conv2d_4_source_30_source_mode <= 5'b0;
      _stream_conv2d_4_source_30_source_offset <= 0;
      _source_stream_conv2d_4_source_30_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_30_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_30_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_30_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_30_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_30_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_30_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_30_pat_stride_3 <= 0;
      _stream_conv2d_4_source_30_source_sel <= 0;
      _stream_conv2d_4_source_30_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_30_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_30_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_30_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_30_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_30_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_30_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_30_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_30_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_30_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_30_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_30_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_30_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_30_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_30_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_30_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_30_pat_stride_buf_3 <= 0;
      __variable_wdata_1837 <= 0;
      _stream_conv2d_4_source_30_source_ram_raddr <= 0;
      _stream_conv2d_4_source_31_source_mode <= 5'b0;
      _stream_conv2d_4_source_31_source_offset <= 0;
      _source_stream_conv2d_4_source_31_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_31_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_31_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_31_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_31_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_31_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_31_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_31_pat_stride_3 <= 0;
      _stream_conv2d_4_source_31_source_sel <= 0;
      _stream_conv2d_4_source_31_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_31_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_31_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_31_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_31_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_31_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_31_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_31_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_31_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_31_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_31_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_31_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_31_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_31_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_31_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_31_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_31_pat_stride_buf_3 <= 0;
      __variable_wdata_1838 <= 0;
      _stream_conv2d_4_source_31_source_ram_raddr <= 0;
      _stream_conv2d_4_source_32_source_mode <= 5'b0;
      _stream_conv2d_4_source_32_source_offset <= 0;
      _source_stream_conv2d_4_source_32_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_32_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_32_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_32_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_32_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_32_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_32_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_32_pat_stride_3 <= 0;
      _stream_conv2d_4_source_32_source_sel <= 0;
      _stream_conv2d_4_source_32_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_32_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_32_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_32_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_32_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_32_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_32_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_32_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_32_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_32_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_32_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_32_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_32_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_32_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_32_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_32_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_32_pat_stride_buf_3 <= 0;
      __variable_wdata_1839 <= 0;
      _stream_conv2d_4_source_32_source_ram_raddr <= 0;
      _stream_conv2d_4_source_33_source_mode <= 5'b0;
      _stream_conv2d_4_source_33_source_offset <= 0;
      _source_stream_conv2d_4_source_33_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_33_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_33_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_33_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_33_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_33_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_33_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_33_pat_stride_3 <= 0;
      _stream_conv2d_4_source_33_source_sel <= 0;
      _stream_conv2d_4_source_33_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_33_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_33_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_33_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_33_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_33_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_33_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_33_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_33_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_33_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_33_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_33_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_33_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_33_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_33_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_33_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_33_pat_stride_buf_3 <= 0;
      __variable_wdata_1840 <= 0;
      _stream_conv2d_4_source_33_source_ram_raddr <= 0;
      _stream_conv2d_4_source_34_source_mode <= 5'b0;
      _stream_conv2d_4_source_34_source_offset <= 0;
      _source_stream_conv2d_4_source_34_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_34_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_34_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_34_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_34_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_34_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_34_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_34_pat_stride_3 <= 0;
      _stream_conv2d_4_source_34_source_sel <= 0;
      _stream_conv2d_4_source_34_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_34_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_34_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_34_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_34_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_34_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_34_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_34_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_34_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_34_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_34_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_34_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_34_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_34_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_34_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_34_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_34_pat_stride_buf_3 <= 0;
      __variable_wdata_1841 <= 0;
      _stream_conv2d_4_source_34_source_ram_raddr <= 0;
      _stream_conv2d_4_source_35_source_mode <= 5'b0;
      _stream_conv2d_4_source_35_source_offset <= 0;
      _source_stream_conv2d_4_source_35_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_35_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_35_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_35_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_35_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_35_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_35_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_35_pat_stride_3 <= 0;
      _stream_conv2d_4_source_35_source_sel <= 0;
      _stream_conv2d_4_source_35_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_35_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_35_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_35_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_35_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_35_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_35_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_35_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_35_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_35_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_35_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_35_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_35_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_35_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_35_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_35_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_35_pat_stride_buf_3 <= 0;
      __variable_wdata_1842 <= 0;
      _stream_conv2d_4_source_35_source_ram_raddr <= 0;
      _stream_conv2d_4_source_36_source_mode <= 5'b0;
      _stream_conv2d_4_source_36_source_offset <= 0;
      _source_stream_conv2d_4_source_36_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_36_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_36_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_36_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_36_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_36_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_36_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_36_pat_stride_3 <= 0;
      _stream_conv2d_4_source_36_source_sel <= 0;
      _stream_conv2d_4_source_36_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_36_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_36_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_36_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_36_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_36_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_36_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_36_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_36_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_36_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_36_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_36_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_36_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_36_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_36_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_36_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_36_pat_stride_buf_3 <= 0;
      __variable_wdata_1843 <= 0;
      _stream_conv2d_4_source_36_source_ram_raddr <= 0;
      _stream_conv2d_4_source_37_source_mode <= 5'b0;
      _stream_conv2d_4_source_37_source_offset <= 0;
      _source_stream_conv2d_4_source_37_pat_size_0 <= 0;
      _source_stream_conv2d_4_source_37_pat_stride_0 <= 0;
      _source_stream_conv2d_4_source_37_pat_size_1 <= 0;
      _source_stream_conv2d_4_source_37_pat_stride_1 <= 0;
      _source_stream_conv2d_4_source_37_pat_size_2 <= 0;
      _source_stream_conv2d_4_source_37_pat_stride_2 <= 0;
      _source_stream_conv2d_4_source_37_pat_size_3 <= 0;
      _source_stream_conv2d_4_source_37_pat_stride_3 <= 0;
      _stream_conv2d_4_source_37_source_sel <= 0;
      _stream_conv2d_4_source_37_source_offset_buf <= 0;
      _source_stream_conv2d_4_source_37_pat_cur_offset_0 <= 0;
      _source_stream_conv2d_4_source_37_pat_cur_offset_1 <= 0;
      _source_stream_conv2d_4_source_37_pat_cur_offset_2 <= 0;
      _source_stream_conv2d_4_source_37_pat_cur_offset_3 <= 0;
      _source_stream_conv2d_4_source_37_pat_count_0 <= 0;
      _source_stream_conv2d_4_source_37_pat_count_1 <= 0;
      _source_stream_conv2d_4_source_37_pat_count_2 <= 0;
      _source_stream_conv2d_4_source_37_pat_count_3 <= 0;
      _source_stream_conv2d_4_source_37_pat_size_buf_0 <= 0;
      _source_stream_conv2d_4_source_37_pat_size_buf_1 <= 0;
      _source_stream_conv2d_4_source_37_pat_size_buf_2 <= 0;
      _source_stream_conv2d_4_source_37_pat_size_buf_3 <= 0;
      _source_stream_conv2d_4_source_37_pat_stride_buf_0 <= 0;
      _source_stream_conv2d_4_source_37_pat_stride_buf_1 <= 0;
      _source_stream_conv2d_4_source_37_pat_stride_buf_2 <= 0;
      _source_stream_conv2d_4_source_37_pat_stride_buf_3 <= 0;
      __variable_wdata_1844 <= 0;
      _stream_conv2d_4_source_37_source_ram_raddr <= 0;
      _tmp_526 <= 0;
      _tmp_527 <= 0;
      _tmp_528 <= 0;
      _tmp_529 <= 0;
      _tmp_530 <= 0;
      _tmp_531 <= 0;
      _tmp_532 <= 0;
      _tmp_533 <= 0;
      _tmp_534 <= 0;
      _tmp_535 <= 0;
      _tmp_536 <= 0;
      _tmp_537 <= 0;
      _tmp_538 <= 0;
      _tmp_539 <= 0;
      _tmp_540 <= 0;
      _tmp_541 <= 0;
      _tmp_542 <= 0;
      _tmp_543 <= 0;
      _tmp_544 <= 0;
      _tmp_545 <= 0;
      _tmp_546 <= 0;
      _tmp_547 <= 0;
      _tmp_548 <= 0;
      _tmp_549 <= 0;
      _tmp_550 <= 0;
      _tmp_551 <= 0;
      _tmp_552 <= 0;
      _tmp_553 <= 0;
      _tmp_554 <= 0;
      _tmp_555 <= 0;
      _tmp_556 <= 0;
      _tmp_557 <= 0;
      _tmp_558 <= 0;
      _tmp_561 <= 0;
      _tmp_562 <= 0;
      _tmp_563 <= 0;
      _tmp_564 <= 0;
      _tmp_565 <= 0;
      _tmp_566 <= 0;
      _tmp_567 <= 0;
      _tmp_568 <= 0;
      _tmp_569 <= 0;
      _tmp_570 <= 0;
      _tmp_571 <= 0;
      _tmp_572 <= 0;
      _tmp_573 <= 0;
      _tmp_574 <= 0;
      _tmp_575 <= 0;
      _tmp_576 <= 0;
      _tmp_577 <= 0;
      _tmp_578 <= 0;
      _tmp_579 <= 0;
      _tmp_580 <= 0;
      _tmp_581 <= 0;
      _tmp_582 <= 0;
      _tmp_583 <= 0;
      _tmp_584 <= 0;
      _tmp_585 <= 0;
      _tmp_586 <= 0;
      _tmp_587 <= 0;
      _tmp_588 <= 0;
      _tmp_589 <= 0;
      _tmp_590 <= 0;
      _tmp_591 <= 0;
      _tmp_592 <= 0;
      _tmp_593 <= 0;
      _tmp_594 <= 0;
      _tmp_595 <= 0;
      _tmp_596 <= 0;
      _tmp_597 <= 0;
      _tmp_598 <= 0;
      _tmp_599 <= 0;
      _tmp_600 <= 0;
      _tmp_601 <= 0;
      _tmp_602 <= 0;
      _tmp_603 <= 0;
      _tmp_604 <= 0;
      _tmp_605 <= 0;
      _tmp_606 <= 0;
      _tmp_607 <= 0;
      _tmp_608 <= 0;
      _tmp_609 <= 0;
      _tmp_610 <= 0;
      _tmp_611 <= 0;
      _tmp_612 <= 0;
      _tmp_613 <= 0;
      _tmp_614 <= 0;
      _tmp_615 <= 0;
      _tmp_616 <= 0;
      _tmp_617 <= 0;
      _tmp_618 <= 0;
      _tmp_619 <= 0;
      _tmp_620 <= 0;
      _tmp_621 <= 0;
      _tmp_622 <= 0;
      _tmp_623 <= 0;
      _tmp_624 <= 0;
      _tmp_625 <= 0;
      _tmp_626 <= 0;
      _stream_conv2d_4_sink_50_sink_mode <= 5'b0;
      _stream_conv2d_4_sink_50_sink_offset <= 0;
      _stream_conv2d_4_sink_50_sink_size <= 0;
      _stream_conv2d_4_sink_50_sink_stride <= 0;
      _stream_conv2d_4_sink_50_sink_sel <= 0;
      _stream_conv2d_4_sink_50_sink_offset_buf <= 0;
      _stream_conv2d_4_sink_50_sink_size_buf <= 0;
      _stream_conv2d_4_sink_50_sink_stride_buf <= 0;
      _stream_conv2d_4_sink_50_sink_waddr <= 0;
      _stream_conv2d_4_sink_50_sink_count <= 0;
      _stream_conv2d_4_sink_50_sink_wdata <= 0;
      _tmp_1017 <= 0;
      _tmp_1018 <= 0;
      _tmp_1019 <= 0;
      _tmp_1020 <= 0;
      _tmp_1021 <= 0;
      _tmp_1022 <= 0;
      __variable_wdata_1553 <= 0;
      _tmp_1023 <= 0;
      _tmp_1024 <= 0;
      _tmp_1025 <= 0;
      _tmp_1026 <= 0;
      _tmp_1029 <= 0;
      _tmp_1032 <= 0;
      _tmp_1033 <= 0;
      _tmp_1034 <= 0;
      _tmp_1035 <= 0;
      _tmp_1036 <= 0;
      _tmp_1037 <= 0;
      _tmp_1038 <= 0;
      _tmp_1039 <= 0;
      _tmp_1040 <= 0;
      _tmp_1041 <= 0;
      _tmp_1042 <= 0;
      _tmp_1043 <= 0;
      _tmp_1044 <= 0;
      _tmp_1045 <= 0;
      _tmp_1046 <= 0;
      _tmp_1047 <= 0;
      _tmp_1048 <= 0;
      _tmp_1049 <= 0;
      _tmp_1050 <= 0;
      _tmp_1051 <= 0;
      _tmp_1052 <= 0;
      _tmp_1053 <= 0;
      _tmp_1054 <= 0;
      _tmp_1055 <= 0;
      _tmp_1056 <= 0;
      _tmp_1057 <= 0;
      _tmp_1058 <= 0;
      _tmp_1059 <= 0;
      _tmp_1060 <= 0;
      _tmp_1061 <= 0;
      _tmp_1062 <= 0;
      _tmp_1063 <= 0;
      _tmp_1064 <= 0;
      _tmp_1065 <= 0;
      _tmp_1066 <= 0;
      _tmp_1067 <= 0;
      _tmp_1068 <= 0;
      _tmp_1069 <= 0;
      _tmp_1070 <= 0;
      _tmp_1071 <= 0;
      _tmp_1072 <= 0;
      _tmp_1073 <= 0;
      _tmp_1074 <= 0;
      _tmp_1075 <= 0;
      _tmp_1076 <= 0;
      _tmp_1077 <= 0;
      _tmp_1078 <= 0;
      _tmp_1079 <= 0;
      _tmp_1080 <= 0;
      _tmp_1081 <= 0;
      _tmp_1082 <= 0;
      _tmp_1083 <= 0;
      _tmp_1084 <= 0;
      _tmp_1085 <= 0;
      _tmp_1086 <= 0;
      _tmp_1087 <= 0;
      _tmp_1088 <= 0;
      _tmp_1089 <= 0;
      _tmp_1090 <= 0;
      _tmp_1091 <= 0;
      _tmp_1092 <= 0;
      _tmp_1093 <= 0;
      _tmp_1094 <= 0;
      _tmp_1095 <= 0;
      _tmp_1096 <= 0;
      _tmp_1097 <= 0;
      _tmp_1098 <= 0;
      _tmp_1099 <= 0;
      _tmp_1100 <= 0;
      _tmp_1101 <= 0;
      _tmp_1102 <= 0;
      _tmp_1103 <= 0;
      _tmp_1104 <= 0;
      _tmp_1105 <= 0;
      _tmp_1106 <= 0;
      _tmp_1107 <= 0;
      _tmp_1108 <= 0;
      _tmp_1109 <= 0;
      _tmp_1110 <= 0;
      _tmp_1111 <= 0;
      _tmp_1112 <= 0;
      _tmp_1113 <= 0;
      _tmp_1114 <= 0;
      _tmp_1115 <= 0;
      _tmp_1116 <= 0;
      _tmp_1117 <= 0;
      _tmp_1118 <= 0;
      _tmp_1119 <= 0;
      _tmp_1120 <= 0;
      _tmp_1121 <= 0;
      _tmp_1122 <= 0;
      _tmp_1123 <= 0;
      _tmp_1124 <= 0;
      _tmp_1125 <= 0;
      _tmp_1126 <= 0;
      _tmp_1127 <= 0;
      _tmp_1128 <= 0;
      _tmp_1129 <= 0;
      _tmp_1130 <= 0;
      _tmp_1131 <= 0;
      _tmp_1132 <= 0;
      _stream_conv2d_4_busy_reg <= 0;
    end else begin
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_7_source_ram_renable <= 0;
        _stream_conv2d_4_source_7_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_7_idle <= _stream_conv2d_4_source_7_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_9_source_ram_renable <= 0;
        _stream_conv2d_4_source_9_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_9_idle <= _stream_conv2d_4_source_9_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_11_source_ram_renable <= 0;
        _stream_conv2d_4_source_11_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_11_idle <= _stream_conv2d_4_source_11_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_13_source_ram_renable <= 0;
        _stream_conv2d_4_source_13_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_13_idle <= _stream_conv2d_4_source_13_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_15_source_ram_renable <= 0;
        _stream_conv2d_4_source_15_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_15_idle <= _stream_conv2d_4_source_15_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_20_source_ram_renable <= 0;
        _stream_conv2d_4_source_20_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_20_idle <= _stream_conv2d_4_source_20_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_21_source_ram_renable <= 0;
        _stream_conv2d_4_source_21_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_21_idle <= _stream_conv2d_4_source_21_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_22_source_ram_renable <= 0;
        _stream_conv2d_4_source_22_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_22_idle <= _stream_conv2d_4_source_22_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_23_source_ram_renable <= 0;
        _stream_conv2d_4_source_23_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_23_idle <= _stream_conv2d_4_source_23_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_24_source_ram_renable <= 0;
        _stream_conv2d_4_source_24_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_24_idle <= _stream_conv2d_4_source_24_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_25_source_ram_renable <= 0;
        _stream_conv2d_4_source_25_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_25_idle <= _stream_conv2d_4_source_25_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_26_source_ram_renable <= 0;
        _stream_conv2d_4_source_26_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_26_idle <= _stream_conv2d_4_source_26_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_27_source_ram_renable <= 0;
        _stream_conv2d_4_source_27_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_27_idle <= _stream_conv2d_4_source_27_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_28_source_ram_renable <= 0;
        _stream_conv2d_4_source_28_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_28_idle <= _stream_conv2d_4_source_28_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_29_source_ram_renable <= 0;
        _stream_conv2d_4_source_29_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_29_idle <= _stream_conv2d_4_source_29_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_30_source_ram_renable <= 0;
        _stream_conv2d_4_source_30_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_30_idle <= _stream_conv2d_4_source_30_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_31_source_ram_renable <= 0;
        _stream_conv2d_4_source_31_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_31_idle <= _stream_conv2d_4_source_31_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_32_source_ram_renable <= 0;
        _stream_conv2d_4_source_32_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_32_idle <= _stream_conv2d_4_source_32_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_33_source_ram_renable <= 0;
        _stream_conv2d_4_source_33_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_33_idle <= _stream_conv2d_4_source_33_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_34_source_ram_renable <= 0;
        _stream_conv2d_4_source_34_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_34_idle <= _stream_conv2d_4_source_34_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_35_source_ram_renable <= 0;
        _stream_conv2d_4_source_35_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_35_idle <= _stream_conv2d_4_source_35_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_36_source_ram_renable <= 0;
        _stream_conv2d_4_source_36_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_36_idle <= _stream_conv2d_4_source_36_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_37_source_ram_renable <= 0;
        _stream_conv2d_4_source_37_source_fifo_deq <= 0;
      end 
      _stream_conv2d_4_source_37_idle <= _stream_conv2d_4_source_37_idle;
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_sink_50_sink_wenable <= 0;
        _stream_conv2d_4_sink_50_sink_fifo_enq <= 0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_sink_51_sink_wenable <= 0;
        _stream_conv2d_4_sink_51_sink_fifo_enq <= 0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_1 <= _stream_conv2d_4_stream_ivalid;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_2 <= __stream_conv2d_4_stream_ivalid_1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_3 <= __stream_conv2d_4_stream_ivalid_2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_4 <= __stream_conv2d_4_stream_ivalid_3;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_5 <= __stream_conv2d_4_stream_ivalid_4;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_6 <= __stream_conv2d_4_stream_ivalid_5;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_7 <= __stream_conv2d_4_stream_ivalid_6;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_8 <= __stream_conv2d_4_stream_ivalid_7;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_9 <= __stream_conv2d_4_stream_ivalid_8;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_10 <= __stream_conv2d_4_stream_ivalid_9;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_11 <= __stream_conv2d_4_stream_ivalid_10;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_12 <= __stream_conv2d_4_stream_ivalid_11;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_13 <= __stream_conv2d_4_stream_ivalid_12;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_14 <= __stream_conv2d_4_stream_ivalid_13;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_15 <= __stream_conv2d_4_stream_ivalid_14;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_16 <= __stream_conv2d_4_stream_ivalid_15;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_17 <= __stream_conv2d_4_stream_ivalid_16;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_18 <= __stream_conv2d_4_stream_ivalid_17;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_19 <= __stream_conv2d_4_stream_ivalid_18;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_20 <= __stream_conv2d_4_stream_ivalid_19;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_21 <= __stream_conv2d_4_stream_ivalid_20;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_22 <= __stream_conv2d_4_stream_ivalid_21;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_23 <= __stream_conv2d_4_stream_ivalid_22;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_24 <= __stream_conv2d_4_stream_ivalid_23;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_25 <= __stream_conv2d_4_stream_ivalid_24;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_26 <= __stream_conv2d_4_stream_ivalid_25;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_27 <= __stream_conv2d_4_stream_ivalid_26;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_28 <= __stream_conv2d_4_stream_ivalid_27;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_29 <= __stream_conv2d_4_stream_ivalid_28;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_30 <= __stream_conv2d_4_stream_ivalid_29;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __stream_conv2d_4_stream_ivalid_31 <= __stream_conv2d_4_stream_ivalid_30;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1611 <= stream_conv2d_4_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1615 <= stream_conv2d_4_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1618 <= stream_conv2d_4_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1621 <= stream_conv2d_4_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1625 <= stream_conv2d_4_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1628 <= stream_conv2d_4_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1631 <= stream_conv2d_4_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1635 <= stream_conv2d_4_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1638 <= stream_conv2d_4_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1641 <= stream_conv2d_4_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1645 <= stream_conv2d_4_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1648 <= stream_conv2d_4_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1651 <= stream_conv2d_4_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1655 <= stream_conv2d_4_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1658 <= stream_conv2d_4_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1661 <= stream_conv2d_4_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1665 <= stream_conv2d_4_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1668 <= stream_conv2d_4_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1671 <= stream_conv2d_4_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1675 <= stream_conv2d_4_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1678 <= stream_conv2d_4_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1681 <= stream_conv2d_4_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1685 <= stream_conv2d_4_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1688 <= stream_conv2d_4_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1691 <= stream_conv2d_4_parameter_1_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1695 <= stream_conv2d_4_parameter_1_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1698 <= stream_conv2d_4_parameter_1_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1701 <= stream_conv2d_4_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1705 <= stream_conv2d_4_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1708 <= stream_conv2d_4_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1711 <= stream_conv2d_4_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1715 <= stream_conv2d_4_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1718 <= stream_conv2d_4_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1721 <= stream_conv2d_4_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1725 <= stream_conv2d_4_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1728 <= stream_conv2d_4_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1731 <= stream_conv2d_4_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1735 <= stream_conv2d_4_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1738 <= stream_conv2d_4_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1741 <= stream_conv2d_4_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1745 <= stream_conv2d_4_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1748 <= stream_conv2d_4_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1751 <= stream_conv2d_4_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1755 <= stream_conv2d_4_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1758 <= stream_conv2d_4_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1761 <= stream_conv2d_4_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1765 <= stream_conv2d_4_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1768 <= stream_conv2d_4_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1771 <= stream_conv2d_4_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1775 <= stream_conv2d_4_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1778 <= stream_conv2d_4_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1781 <= stream_conv2d_4_parameter_2_data == 3'sd2;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1785 <= stream_conv2d_4_parameter_2_data == 2'sd1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _eq_data_1788 <= stream_conv2d_4_parameter_2_data == 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_1943 <= _cond_data_1583 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_1962 <= _cond_data_1583 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_1981 <= _cond_data_1583 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_2000 <= _cond_data_1583 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_2019 <= _cond_data_1583 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_2038 <= _cond_data_1583 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_2057 <= _cond_data_1583 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_2076 <= _cond_data_1583 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_2095 <= _cond_data_1583 + stream_conv2d_4_parameter_16_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_2111 <= _cond_data_1590 + stream_conv2d_4_parameter_17_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_2130 <= _cond_data_1597 + stream_conv2d_4_parameter_18_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2258__variable_1604 <= stream_conv2d_4_source_22_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2259__variable_1603 <= stream_conv2d_4_source_21_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2260__variable_1602 <= stream_conv2d_4_source_20_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2261__variable_1607 <= stream_conv2d_4_source_25_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2262__variable_1606 <= stream_conv2d_4_source_24_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2263__variable_1605 <= stream_conv2d_4_source_23_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2264__variable_1610 <= stream_conv2d_4_source_28_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2265__variable_1609 <= stream_conv2d_4_source_27_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2266__variable_1608 <= stream_conv2d_4_source_26_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2267_pointer_1890 <= _pointer_data_1890;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2268_reinterpretcast_1881 <= _reinterpretcast_data_1881;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2269_pointer_1892 <= _pointer_data_1892;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2270_reinterpretcast_1882 <= _reinterpretcast_data_1882;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2271_pointer_1894 <= _pointer_data_1894;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2272_reinterpretcast_1883 <= _reinterpretcast_data_1883;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2273_pointer_1896 <= _pointer_data_1896;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2274_reinterpretcast_1884 <= _reinterpretcast_data_1884;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2275_pointer_1898 <= _pointer_data_1898;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2276_reinterpretcast_1885 <= _reinterpretcast_data_1885;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2277_pointer_1900 <= _pointer_data_1900;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2278_reinterpretcast_1886 <= _reinterpretcast_data_1886;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2279_pointer_1902 <= _pointer_data_1902;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2280_reinterpretcast_1887 <= _reinterpretcast_data_1887;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2281_pointer_1904 <= _pointer_data_1904;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2282_reinterpretcast_1888 <= _reinterpretcast_data_1888;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2283_pointer_1906 <= _pointer_data_1906;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2284_reinterpretcast_1889 <= _reinterpretcast_data_1889;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2285__variable_1553 <= stream_conv2d_4__reduce_reset_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2310__variable_1548 <= stream_conv2d_4_parameter_0_data;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2323_cond_1569 <= _cond_data_1569;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2342_cond_1576 <= _cond_data_1576;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2286__delay_2285__variable_1553 <= __delay_data_2285__variable_1553;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2298_plus_2111 <= _plus_data_2111;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2311__delay_2310__variable_1548 <= __delay_data_2310__variable_1548;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2324__delay_2323_cond_1569 <= __delay_data_2323_cond_1569;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2343__delay_2342_cond_1576 <= __delay_data_2342_cond_1576;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2362_plus_2130 <= _plus_data_2130;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2287__delay_2286__delay_2285__variable_1553 <= __delay_data_2286__delay_2285__variable_1553;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2299__delay_2298_plus_2111 <= __delay_data_2298_plus_2111;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2312__delay_2311__delay_2310__variable_1548 <= __delay_data_2311__delay_2310__variable_1548;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2325__delay_2324__delay_2323_cond_1569 <= __delay_data_2324__delay_2323_cond_1569;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2344__delay_2343__delay_2342_cond_1576 <= __delay_data_2343__delay_2342_cond_1576;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2363__delay_2362_plus_2130 <= __delay_data_2362_plus_2130;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2288__delay_2287__delay_2286____variable_1553 <= __delay_data_2287__delay_2286__delay_2285__variable_1553;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2300__delay_2299__delay_2298_plus_2111 <= __delay_data_2299__delay_2298_plus_2111;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2313__delay_2312__delay_2311____variable_1548 <= __delay_data_2312__delay_2311__delay_2310__variable_1548;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2326__delay_2325__delay_2324___cond_1569 <= __delay_data_2325__delay_2324__delay_2323_cond_1569;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2345__delay_2344__delay_2343___cond_1576 <= __delay_data_2344__delay_2343__delay_2342_cond_1576;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2364__delay_2363__delay_2362_plus_2130 <= __delay_data_2363__delay_2362_plus_2130;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2289__delay_2288__delay_2287____variable_1553 <= __delay_data_2288__delay_2287__delay_2286____variable_1553;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2301__delay_2300__delay_2299___plus_2111 <= __delay_data_2300__delay_2299__delay_2298_plus_2111;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2314__delay_2313__delay_2312____variable_1548 <= __delay_data_2313__delay_2312__delay_2311____variable_1548;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2327__delay_2326__delay_2325___cond_1569 <= __delay_data_2326__delay_2325__delay_2324___cond_1569;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2346__delay_2345__delay_2344___cond_1576 <= __delay_data_2345__delay_2344__delay_2343___cond_1576;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2365__delay_2364__delay_2363___plus_2130 <= __delay_data_2364__delay_2363__delay_2362_plus_2130;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2290__delay_2289__delay_2288____variable_1553 <= __delay_data_2289__delay_2288__delay_2287____variable_1553;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2302__delay_2301__delay_2300___plus_2111 <= __delay_data_2301__delay_2300__delay_2299___plus_2111;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2315__delay_2314__delay_2313____variable_1548 <= __delay_data_2314__delay_2313__delay_2312____variable_1548;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2328__delay_2327__delay_2326___cond_1569 <= __delay_data_2327__delay_2326__delay_2325___cond_1569;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2347__delay_2346__delay_2345___cond_1576 <= __delay_data_2346__delay_2345__delay_2344___cond_1576;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2366__delay_2365__delay_2364___plus_2130 <= __delay_data_2365__delay_2364__delay_2363___plus_2130;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2291__delay_2290__delay_2289____variable_1553 <= __delay_data_2290__delay_2289__delay_2288____variable_1553;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2303__delay_2302__delay_2301___plus_2111 <= __delay_data_2302__delay_2301__delay_2300___plus_2111;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2316__delay_2315__delay_2314____variable_1548 <= __delay_data_2315__delay_2314__delay_2313____variable_1548;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2329__delay_2328__delay_2327___cond_1569 <= __delay_data_2328__delay_2327__delay_2326___cond_1569;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2348__delay_2347__delay_2346___cond_1576 <= __delay_data_2347__delay_2346__delay_2345___cond_1576;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2367__delay_2366__delay_2365___plus_2130 <= __delay_data_2366__delay_2365__delay_2364___plus_2130;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2292__delay_2291__delay_2290____variable_1553 <= __delay_data_2291__delay_2290__delay_2289____variable_1553;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2304__delay_2303__delay_2302___plus_2111 <= __delay_data_2303__delay_2302__delay_2301___plus_2111;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2317__delay_2316__delay_2315____variable_1548 <= __delay_data_2316__delay_2315__delay_2314____variable_1548;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2330__delay_2329__delay_2328___cond_1569 <= __delay_data_2329__delay_2328__delay_2327___cond_1569;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2349__delay_2348__delay_2347___cond_1576 <= __delay_data_2348__delay_2347__delay_2346___cond_1576;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2368__delay_2367__delay_2366___plus_2130 <= __delay_data_2367__delay_2366__delay_2365___plus_2130;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2293__delay_2292__delay_2291____variable_1553 <= __delay_data_2292__delay_2291__delay_2290____variable_1553;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2305__delay_2304__delay_2303___plus_2111 <= __delay_data_2304__delay_2303__delay_2302___plus_2111;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2318__delay_2317__delay_2316____variable_1548 <= __delay_data_2317__delay_2316__delay_2315____variable_1548;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2331__delay_2330__delay_2329___cond_1569 <= __delay_data_2330__delay_2329__delay_2328___cond_1569;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2350__delay_2349__delay_2348___cond_1576 <= __delay_data_2349__delay_2348__delay_2347___cond_1576;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2369__delay_2368__delay_2367___plus_2130 <= __delay_data_2368__delay_2367__delay_2366___plus_2130;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2294__delay_2293__delay_2292____variable_1553 <= __delay_data_2293__delay_2292__delay_2291____variable_1553;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2306__delay_2305__delay_2304___plus_2111 <= __delay_data_2305__delay_2304__delay_2303___plus_2111;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2319__delay_2318__delay_2317____variable_1548 <= __delay_data_2318__delay_2317__delay_2316____variable_1548;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2332__delay_2331__delay_2330___cond_1569 <= __delay_data_2331__delay_2330__delay_2329___cond_1569;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2351__delay_2350__delay_2349___cond_1576 <= __delay_data_2350__delay_2349__delay_2348___cond_1576;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2370__delay_2369__delay_2368___plus_2130 <= __delay_data_2369__delay_2368__delay_2367___plus_2130;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2295__delay_2294__delay_2293____variable_1553 <= __delay_data_2294__delay_2293__delay_2292____variable_1553;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2307__delay_2306__delay_2305___plus_2111 <= __delay_data_2306__delay_2305__delay_2304___plus_2111;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2320__delay_2319__delay_2318____variable_1548 <= __delay_data_2319__delay_2318__delay_2317____variable_1548;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2333__delay_2332__delay_2331___cond_1569 <= __delay_data_2332__delay_2331__delay_2330___cond_1569;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2352__delay_2351__delay_2350___cond_1576 <= __delay_data_2351__delay_2350__delay_2349___cond_1576;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2371__delay_2370__delay_2369___plus_2130 <= __delay_data_2370__delay_2369__delay_2368___plus_2130;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2296__delay_2295__delay_2294____variable_1553 <= __delay_data_2295__delay_2294__delay_2293____variable_1553;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2308__delay_2307__delay_2306___plus_2111 <= __delay_data_2307__delay_2306__delay_2305___plus_2111;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2321__delay_2320__delay_2319____variable_1548 <= __delay_data_2320__delay_2319__delay_2318____variable_1548;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2334__delay_2333__delay_2332___cond_1569 <= __delay_data_2333__delay_2332__delay_2331___cond_1569;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2353__delay_2352__delay_2351___cond_1576 <= __delay_data_2352__delay_2351__delay_2350___cond_1576;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2372__delay_2371__delay_2370___plus_2130 <= __delay_data_2371__delay_2370__delay_2369___plus_2130;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2297__delay_2296__delay_2295____variable_1553 <= __delay_data_2296__delay_2295__delay_2294____variable_1553;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2309__delay_2308__delay_2307___plus_2111 <= __delay_data_2308__delay_2307__delay_2306___plus_2111;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2322__delay_2321__delay_2320____variable_1548 <= __delay_data_2321__delay_2320__delay_2319____variable_1548;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2335__delay_2334__delay_2333___cond_1569 <= __delay_data_2334__delay_2333__delay_2332___cond_1569;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2354__delay_2353__delay_2352___cond_1576 <= __delay_data_2353__delay_2352__delay_2351___cond_1576;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2373__delay_2372__delay_2371___plus_2130 <= __delay_data_2372__delay_2371__delay_2370___plus_2130;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2336__delay_2335__delay_2334___cond_1569 <= __delay_data_2335__delay_2334__delay_2333___cond_1569;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2355__delay_2354__delay_2353___cond_1576 <= __delay_data_2354__delay_2353__delay_2352___cond_1576;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2374__delay_2373__delay_2372___plus_2130 <= __delay_data_2373__delay_2372__delay_2371___plus_2130;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2337__delay_2336__delay_2335___cond_1569 <= __delay_data_2336__delay_2335__delay_2334___cond_1569;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2356__delay_2355__delay_2354___cond_1576 <= __delay_data_2355__delay_2354__delay_2353___cond_1576;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2375__delay_2374__delay_2373___plus_2130 <= __delay_data_2374__delay_2373__delay_2372___plus_2130;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2338__delay_2337__delay_2336___cond_1569 <= __delay_data_2337__delay_2336__delay_2335___cond_1569;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2357__delay_2356__delay_2355___cond_1576 <= __delay_data_2356__delay_2355__delay_2354___cond_1576;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2376__delay_2375__delay_2374___plus_2130 <= __delay_data_2375__delay_2374__delay_2373___plus_2130;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2339__delay_2338__delay_2337___cond_1569 <= __delay_data_2338__delay_2337__delay_2336___cond_1569;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2358__delay_2357__delay_2356___cond_1576 <= __delay_data_2357__delay_2356__delay_2355___cond_1576;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2377__delay_2376__delay_2375___plus_2130 <= __delay_data_2376__delay_2375__delay_2374___plus_2130;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2340__delay_2339__delay_2338___cond_1569 <= __delay_data_2339__delay_2338__delay_2337___cond_1569;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2359__delay_2358__delay_2357___cond_1576 <= __delay_data_2358__delay_2357__delay_2356___cond_1576;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2378__delay_2377__delay_2376___plus_2130 <= __delay_data_2377__delay_2376__delay_2375___plus_2130;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2341__delay_2340__delay_2339___cond_1569 <= __delay_data_2340__delay_2339__delay_2338___cond_1569;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2360__delay_2359__delay_2358___cond_1576 <= __delay_data_2359__delay_2358__delay_2357___cond_1576;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2379__delay_2378__delay_2377___plus_2130 <= __delay_data_2378__delay_2377__delay_2376___plus_2130;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _plus_data_2114 <= __substreamoutput_data_2112 + __delay_data_2341__delay_2340__delay_2339___cond_1569;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2361__delay_2360__delay_2359___cond_1576 <= __delay_data_2360__delay_2359__delay_2358___cond_1576;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2380__delay_2379__delay_2378___plus_2130 <= __delay_data_2379__delay_2378__delay_2377___plus_2130;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2382__substreamoutput_2113 <= __substreamoutput_data_2113;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2383__delay_2382__substreamoutput_2113 <= __delay_data_2382__substreamoutput_2113;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2384__delay_2383____substreamoutput_2113 <= __delay_data_2383__delay_2382__substreamoutput_2113;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2385__delay_2384____substreamoutput_2113 <= __delay_data_2384__delay_2383____substreamoutput_2113;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2386__delay_2385____substreamoutput_2113 <= __delay_data_2385__delay_2384____substreamoutput_2113;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2387__delay_2386____substreamoutput_2113 <= __delay_data_2386__delay_2385____substreamoutput_2113;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2388__delay_2387____substreamoutput_2113 <= __delay_data_2387__delay_2386____substreamoutput_2113;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2389__delay_2388____substreamoutput_2113 <= __delay_data_2388__delay_2387____substreamoutput_2113;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2390__delay_2389____substreamoutput_2113 <= __delay_data_2389__delay_2388____substreamoutput_2113;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2391__delay_2390____substreamoutput_2113 <= __delay_data_2390__delay_2389____substreamoutput_2113;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _greaterthan_data_2133 <= __substreamoutput_data_2131 > 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2381__substreamoutput_2131 <= __substreamoutput_data_2131;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2392__delay_2391____substreamoutput_2113 <= __delay_data_2391__delay_2390____substreamoutput_2113;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _cond_data_2135 <= (_greaterthan_data_2133)? __delay_data_2381__substreamoutput_2131 : 1'sd0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        __delay_data_2393__delay_2392____substreamoutput_2113 <= __delay_data_2392__delay_2391____substreamoutput_2113;
      end 
      if(_set_flag_328) begin
        _stream_conv2d_4_parameter_0_next_parameter_data <= cparam_conv2d_4_stream_reduce_size;
      end 
      if(_stream_conv2d_4_source_start) begin
        __variable_wdata_1548 <= _stream_conv2d_4_parameter_0_next_parameter_data;
      end 
      if(_set_flag_329) begin
        _stream_conv2d_4_parameter_1_next_parameter_data <= conv2d_4_col_select;
      end 
      if(_stream_conv2d_4_source_start) begin
        __variable_wdata_1549 <= _stream_conv2d_4_parameter_1_next_parameter_data;
      end 
      if(_set_flag_330) begin
        _stream_conv2d_4_parameter_2_next_parameter_data <= conv2d_4_row_select_buf;
      end 
      if(_stream_conv2d_4_source_start) begin
        __variable_wdata_1550 <= _stream_conv2d_4_parameter_2_next_parameter_data;
      end 
      if(_set_flag_331) begin
        _stream_conv2d_4_parameter_3_next_parameter_data <= conv2d_4_stream_pad_masks;
      end 
      if(_stream_conv2d_4_source_start) begin
        __variable_wdata_1551 <= _stream_conv2d_4_parameter_3_next_parameter_data;
      end 
      if(_set_flag_332) begin
        _stream_conv2d_4_parameter_4_next_parameter_data <= cparam_conv2d_4_stream_omit_mask;
      end 
      if(_stream_conv2d_4_source_start) begin
        __variable_wdata_1552 <= _stream_conv2d_4_parameter_4_next_parameter_data;
      end 
      if(_set_flag_333) begin
        _stream_conv2d_4_parameter_6_next_parameter_data <= cparam_conv2d_4_bias_scala;
      end 
      if(_stream_conv2d_4_source_start) begin
        __variable_wdata_1563 <= _stream_conv2d_4_parameter_6_next_parameter_data;
      end 
      if(_set_flag_334) begin
        _stream_conv2d_4_source_7_source_mode <= 5'b10;
        _stream_conv2d_4_source_7_source_offset <= (cparam_conv2d_4_bias_num == 1)? 0 : conv2d_4_och_count_buf;
      end 
      if(_set_flag_334) begin
        _source_stream_conv2d_4_source_7_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_7_pat_stride_0 <= 0;
      end 
      if(_set_flag_334) begin
        _source_stream_conv2d_4_source_7_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_7_pat_stride_1 <= (cparam_conv2d_4_bias_num == 1)? 0 : 1;
      end 
      if(_set_flag_334) begin
        _source_stream_conv2d_4_source_7_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_7_pat_stride_2 <= 0;
      end 
      if(_set_flag_334) begin
        _source_stream_conv2d_4_source_7_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_7_pat_stride_3 <= 0;
      end 
      if(_set_flag_334) begin
        _stream_conv2d_4_source_7_source_sel <= 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_7_source_offset_buf <= _stream_conv2d_4_source_7_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_count_0 <= _source_stream_conv2d_4_source_7_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_count_1 <= _source_stream_conv2d_4_source_7_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_count_2 <= _source_stream_conv2d_4_source_7_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_count_3 <= _source_stream_conv2d_4_source_7_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_size_buf_0 <= _source_stream_conv2d_4_source_7_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_size_buf_1 <= _source_stream_conv2d_4_source_7_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_size_buf_2 <= _source_stream_conv2d_4_source_7_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_size_buf_3 <= _source_stream_conv2d_4_source_7_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_stride_buf_0 <= _source_stream_conv2d_4_source_7_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_stride_buf_1 <= _source_stream_conv2d_4_source_7_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_stride_buf_2 <= _source_stream_conv2d_4_source_7_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_stride_buf_3 <= _source_stream_conv2d_4_source_7_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_1564 <= _stream_conv2d_4_source_7_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_7_source_pat_fsm_0 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_7_idle <= 0;
        _stream_conv2d_4_source_7_source_ram_raddr <= _stream_conv2d_4_source_7_source_pat_all_offset;
        _stream_conv2d_4_source_7_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_7_source_pat_fsm_0 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_cur_offset_0 <= _source_stream_conv2d_4_source_7_pat_cur_offset_0 + _source_stream_conv2d_4_source_7_pat_stride_buf_0;
        _source_stream_conv2d_4_source_7_pat_count_0 <= _source_stream_conv2d_4_source_7_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_7_source_pat_fsm_0 == 1) && (_source_stream_conv2d_4_source_7_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_7_pat_count_0 <= _source_stream_conv2d_4_source_7_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_7_source_pat_fsm_0 == 1) && (_source_stream_conv2d_4_source_7_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_cur_offset_1 <= _source_stream_conv2d_4_source_7_pat_cur_offset_1 + _source_stream_conv2d_4_source_7_pat_stride_buf_1;
        _source_stream_conv2d_4_source_7_pat_count_1 <= _source_stream_conv2d_4_source_7_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_7_source_pat_fsm_0 == 1) && (_source_stream_conv2d_4_source_7_pat_count_0 == 0) && (_source_stream_conv2d_4_source_7_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_7_pat_count_1 <= _source_stream_conv2d_4_source_7_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_7_source_pat_fsm_0 == 1) && ((_source_stream_conv2d_4_source_7_pat_count_0 == 0) && (_source_stream_conv2d_4_source_7_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_cur_offset_2 <= _source_stream_conv2d_4_source_7_pat_cur_offset_2 + _source_stream_conv2d_4_source_7_pat_stride_buf_2;
        _source_stream_conv2d_4_source_7_pat_count_2 <= _source_stream_conv2d_4_source_7_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_7_source_pat_fsm_0 == 1) && ((_source_stream_conv2d_4_source_7_pat_count_0 == 0) && (_source_stream_conv2d_4_source_7_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_7_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_7_pat_count_2 <= _source_stream_conv2d_4_source_7_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_7_source_pat_fsm_0 == 1) && ((_source_stream_conv2d_4_source_7_pat_count_0 == 0) && (_source_stream_conv2d_4_source_7_pat_count_1 == 0) && (_source_stream_conv2d_4_source_7_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_cur_offset_3 <= _source_stream_conv2d_4_source_7_pat_cur_offset_3 + _source_stream_conv2d_4_source_7_pat_stride_buf_3;
        _source_stream_conv2d_4_source_7_pat_count_3 <= _source_stream_conv2d_4_source_7_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_7_source_pat_fsm_0 == 1) && ((_source_stream_conv2d_4_source_7_pat_count_0 == 0) && (_source_stream_conv2d_4_source_7_pat_count_1 == 0) && (_source_stream_conv2d_4_source_7_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_7_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_7_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_7_pat_count_3 <= _source_stream_conv2d_4_source_7_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_7_source_pat_fsm_0 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_7_source_ram_renable <= 0;
        _stream_conv2d_4_source_7_idle <= 1;
      end 
      if((_stream_conv2d_4_source_7_source_pat_fsm_0 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_7_source_ram_renable <= 0;
        _stream_conv2d_4_source_7_idle <= 1;
      end 
      if(_set_flag_343) begin
        _stream_conv2d_4_parameter_8_next_parameter_data <= cparam_conv2d_4_scale_scala;
      end 
      if(_stream_conv2d_4_source_start) begin
        __variable_wdata_1570 <= _stream_conv2d_4_parameter_8_next_parameter_data;
      end 
      if(_set_flag_344) begin
        _stream_conv2d_4_source_9_source_mode <= 5'b10;
        _stream_conv2d_4_source_9_source_offset <= (cparam_conv2d_4_scale_num == 1)? 0 : conv2d_4_och_count_buf;
      end 
      if(_set_flag_344) begin
        _source_stream_conv2d_4_source_9_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_9_pat_stride_0 <= 0;
      end 
      if(_set_flag_344) begin
        _source_stream_conv2d_4_source_9_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_9_pat_stride_1 <= (cparam_conv2d_4_scale_num == 1)? 0 : 1;
      end 
      if(_set_flag_344) begin
        _source_stream_conv2d_4_source_9_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_9_pat_stride_2 <= 0;
      end 
      if(_set_flag_344) begin
        _source_stream_conv2d_4_source_9_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_9_pat_stride_3 <= 0;
      end 
      if(_set_flag_344) begin
        _stream_conv2d_4_source_9_source_sel <= 2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_9_source_offset_buf <= _stream_conv2d_4_source_9_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_count_0 <= _source_stream_conv2d_4_source_9_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_count_1 <= _source_stream_conv2d_4_source_9_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_count_2 <= _source_stream_conv2d_4_source_9_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_count_3 <= _source_stream_conv2d_4_source_9_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_size_buf_0 <= _source_stream_conv2d_4_source_9_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_size_buf_1 <= _source_stream_conv2d_4_source_9_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_size_buf_2 <= _source_stream_conv2d_4_source_9_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_size_buf_3 <= _source_stream_conv2d_4_source_9_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_stride_buf_0 <= _source_stream_conv2d_4_source_9_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_stride_buf_1 <= _source_stream_conv2d_4_source_9_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_stride_buf_2 <= _source_stream_conv2d_4_source_9_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_stride_buf_3 <= _source_stream_conv2d_4_source_9_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_1571 <= _stream_conv2d_4_source_9_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_9_source_pat_fsm_1 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_9_idle <= 0;
        _stream_conv2d_4_source_9_source_ram_raddr <= _stream_conv2d_4_source_9_source_pat_all_offset;
        _stream_conv2d_4_source_9_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_9_source_pat_fsm_1 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_cur_offset_0 <= _source_stream_conv2d_4_source_9_pat_cur_offset_0 + _source_stream_conv2d_4_source_9_pat_stride_buf_0;
        _source_stream_conv2d_4_source_9_pat_count_0 <= _source_stream_conv2d_4_source_9_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_9_source_pat_fsm_1 == 1) && (_source_stream_conv2d_4_source_9_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_9_pat_count_0 <= _source_stream_conv2d_4_source_9_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_9_source_pat_fsm_1 == 1) && (_source_stream_conv2d_4_source_9_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_cur_offset_1 <= _source_stream_conv2d_4_source_9_pat_cur_offset_1 + _source_stream_conv2d_4_source_9_pat_stride_buf_1;
        _source_stream_conv2d_4_source_9_pat_count_1 <= _source_stream_conv2d_4_source_9_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_9_source_pat_fsm_1 == 1) && (_source_stream_conv2d_4_source_9_pat_count_0 == 0) && (_source_stream_conv2d_4_source_9_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_9_pat_count_1 <= _source_stream_conv2d_4_source_9_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_9_source_pat_fsm_1 == 1) && ((_source_stream_conv2d_4_source_9_pat_count_0 == 0) && (_source_stream_conv2d_4_source_9_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_cur_offset_2 <= _source_stream_conv2d_4_source_9_pat_cur_offset_2 + _source_stream_conv2d_4_source_9_pat_stride_buf_2;
        _source_stream_conv2d_4_source_9_pat_count_2 <= _source_stream_conv2d_4_source_9_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_9_source_pat_fsm_1 == 1) && ((_source_stream_conv2d_4_source_9_pat_count_0 == 0) && (_source_stream_conv2d_4_source_9_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_9_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_9_pat_count_2 <= _source_stream_conv2d_4_source_9_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_9_source_pat_fsm_1 == 1) && ((_source_stream_conv2d_4_source_9_pat_count_0 == 0) && (_source_stream_conv2d_4_source_9_pat_count_1 == 0) && (_source_stream_conv2d_4_source_9_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_cur_offset_3 <= _source_stream_conv2d_4_source_9_pat_cur_offset_3 + _source_stream_conv2d_4_source_9_pat_stride_buf_3;
        _source_stream_conv2d_4_source_9_pat_count_3 <= _source_stream_conv2d_4_source_9_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_9_source_pat_fsm_1 == 1) && ((_source_stream_conv2d_4_source_9_pat_count_0 == 0) && (_source_stream_conv2d_4_source_9_pat_count_1 == 0) && (_source_stream_conv2d_4_source_9_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_9_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_9_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_9_pat_count_3 <= _source_stream_conv2d_4_source_9_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_9_source_pat_fsm_1 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_9_source_ram_renable <= 0;
        _stream_conv2d_4_source_9_idle <= 1;
      end 
      if((_stream_conv2d_4_source_9_source_pat_fsm_1 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_9_source_ram_renable <= 0;
        _stream_conv2d_4_source_9_idle <= 1;
      end 
      if(_set_flag_353) begin
        _stream_conv2d_4_parameter_10_next_parameter_data <= 1;
      end 
      if(_stream_conv2d_4_source_start) begin
        __variable_wdata_1577 <= _stream_conv2d_4_parameter_10_next_parameter_data;
      end 
      if(_set_flag_354) begin
        _stream_conv2d_4_source_11_source_mode <= 5'b0;
        _stream_conv2d_4_source_11_source_empty_data <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_stream_oready && !(|(_stream_conv2d_4_source_11_source_mode & 5'b0))) begin
        _stream_conv2d_4_source_11_idle <= 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_stream_oready && !(|(_stream_conv2d_4_source_11_source_mode & 5'b0)) && _stream_conv2d_4_is_root) begin
        __variable_wdata_1578 <= _stream_conv2d_4_source_11_source_empty_data;
      end 
      if(_set_flag_355) begin
        _stream_conv2d_4_parameter_12_next_parameter_data <= 1;
      end 
      if(_stream_conv2d_4_source_start) begin
        __variable_wdata_1584 <= _stream_conv2d_4_parameter_12_next_parameter_data;
      end 
      if(_set_flag_356) begin
        _stream_conv2d_4_source_13_source_mode <= 5'b0;
        _stream_conv2d_4_source_13_source_empty_data <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_stream_oready && !(|(_stream_conv2d_4_source_13_source_mode & 5'b0))) begin
        _stream_conv2d_4_source_13_idle <= 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_stream_oready && !(|(_stream_conv2d_4_source_13_source_mode & 5'b0)) && _stream_conv2d_4_is_root) begin
        __variable_wdata_1585 <= _stream_conv2d_4_source_13_source_empty_data;
      end 
      if(_set_flag_357) begin
        _stream_conv2d_4_parameter_14_next_parameter_data <= 1;
      end 
      if(_stream_conv2d_4_source_start) begin
        __variable_wdata_1591 <= _stream_conv2d_4_parameter_14_next_parameter_data;
      end 
      if(_set_flag_358) begin
        _stream_conv2d_4_source_15_source_mode <= 5'b0;
        _stream_conv2d_4_source_15_source_empty_data <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_stream_oready && !(|(_stream_conv2d_4_source_15_source_mode & 5'b0))) begin
        _stream_conv2d_4_source_15_idle <= 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_stream_oready && !(|(_stream_conv2d_4_source_15_source_mode & 5'b0)) && _stream_conv2d_4_is_root) begin
        __variable_wdata_1592 <= _stream_conv2d_4_source_15_source_empty_data;
      end 
      if(_set_flag_359) begin
        _stream_conv2d_4_parameter_16_next_parameter_data <= cparam_conv2d_4_cshamt_mul_value;
      end 
      if(_stream_conv2d_4_source_start) begin
        __variable_wdata_1598 <= _stream_conv2d_4_parameter_16_next_parameter_data;
      end 
      if(_set_flag_360) begin
        _stream_conv2d_4_parameter_17_next_parameter_data <= cparam_conv2d_4_cshamt_sum_value;
      end 
      if(_stream_conv2d_4_source_start) begin
        __variable_wdata_1599 <= _stream_conv2d_4_parameter_17_next_parameter_data;
      end 
      if(_set_flag_361) begin
        _stream_conv2d_4_parameter_18_next_parameter_data <= cparam_conv2d_4_cshamt_out_value;
      end 
      if(_stream_conv2d_4_source_start) begin
        __variable_wdata_1600 <= _stream_conv2d_4_parameter_18_next_parameter_data;
      end 
      if(_set_flag_362) begin
        _stream_conv2d_4_parameter_19_next_parameter_data <= cparam_conv2d_4_act_func_index;
      end 
      if(_stream_conv2d_4_source_start) begin
        __variable_wdata_1601 <= _stream_conv2d_4_parameter_19_next_parameter_data;
      end 
      if(_set_flag_363) begin
        _stream_conv2d_4_source_20_source_mode <= 5'b10;
        _stream_conv2d_4_source_20_source_offset <= conv2d_4_stream_act_local_0 + conv2d_4_act_page_comp_offset_buf_0;
      end 
      if(_set_flag_363) begin
        _source_stream_conv2d_4_source_20_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_20_pat_stride_0 <= 1;
      end 
      if(_set_flag_363) begin
        _source_stream_conv2d_4_source_20_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_20_pat_stride_1 <= 0;
      end 
      if(_set_flag_363) begin
        _source_stream_conv2d_4_source_20_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_20_pat_stride_2 <= 0;
      end 
      if(_set_flag_363) begin
        _source_stream_conv2d_4_source_20_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_20_pat_stride_3 <= 0;
      end 
      if(_set_flag_363) begin
        _stream_conv2d_4_source_20_source_sel <= 3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_20_source_offset_buf <= _stream_conv2d_4_source_20_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_count_0 <= _source_stream_conv2d_4_source_20_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_count_1 <= _source_stream_conv2d_4_source_20_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_count_2 <= _source_stream_conv2d_4_source_20_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_count_3 <= _source_stream_conv2d_4_source_20_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_size_buf_0 <= _source_stream_conv2d_4_source_20_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_size_buf_1 <= _source_stream_conv2d_4_source_20_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_size_buf_2 <= _source_stream_conv2d_4_source_20_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_size_buf_3 <= _source_stream_conv2d_4_source_20_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_stride_buf_0 <= _source_stream_conv2d_4_source_20_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_stride_buf_1 <= _source_stream_conv2d_4_source_20_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_stride_buf_2 <= _source_stream_conv2d_4_source_20_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_stride_buf_3 <= _source_stream_conv2d_4_source_20_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_1602 <= _stream_conv2d_4_source_20_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_20_source_pat_fsm_2 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_20_idle <= 0;
        _stream_conv2d_4_source_20_source_ram_raddr <= _stream_conv2d_4_source_20_source_pat_all_offset;
        _stream_conv2d_4_source_20_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_20_source_pat_fsm_2 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_cur_offset_0 <= _source_stream_conv2d_4_source_20_pat_cur_offset_0 + _source_stream_conv2d_4_source_20_pat_stride_buf_0;
        _source_stream_conv2d_4_source_20_pat_count_0 <= _source_stream_conv2d_4_source_20_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_20_source_pat_fsm_2 == 1) && (_source_stream_conv2d_4_source_20_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_20_pat_count_0 <= _source_stream_conv2d_4_source_20_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_20_source_pat_fsm_2 == 1) && (_source_stream_conv2d_4_source_20_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_cur_offset_1 <= _source_stream_conv2d_4_source_20_pat_cur_offset_1 + _source_stream_conv2d_4_source_20_pat_stride_buf_1;
        _source_stream_conv2d_4_source_20_pat_count_1 <= _source_stream_conv2d_4_source_20_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_20_source_pat_fsm_2 == 1) && (_source_stream_conv2d_4_source_20_pat_count_0 == 0) && (_source_stream_conv2d_4_source_20_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_20_pat_count_1 <= _source_stream_conv2d_4_source_20_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_20_source_pat_fsm_2 == 1) && ((_source_stream_conv2d_4_source_20_pat_count_0 == 0) && (_source_stream_conv2d_4_source_20_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_cur_offset_2 <= _source_stream_conv2d_4_source_20_pat_cur_offset_2 + _source_stream_conv2d_4_source_20_pat_stride_buf_2;
        _source_stream_conv2d_4_source_20_pat_count_2 <= _source_stream_conv2d_4_source_20_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_20_source_pat_fsm_2 == 1) && ((_source_stream_conv2d_4_source_20_pat_count_0 == 0) && (_source_stream_conv2d_4_source_20_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_20_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_20_pat_count_2 <= _source_stream_conv2d_4_source_20_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_20_source_pat_fsm_2 == 1) && ((_source_stream_conv2d_4_source_20_pat_count_0 == 0) && (_source_stream_conv2d_4_source_20_pat_count_1 == 0) && (_source_stream_conv2d_4_source_20_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_cur_offset_3 <= _source_stream_conv2d_4_source_20_pat_cur_offset_3 + _source_stream_conv2d_4_source_20_pat_stride_buf_3;
        _source_stream_conv2d_4_source_20_pat_count_3 <= _source_stream_conv2d_4_source_20_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_20_source_pat_fsm_2 == 1) && ((_source_stream_conv2d_4_source_20_pat_count_0 == 0) && (_source_stream_conv2d_4_source_20_pat_count_1 == 0) && (_source_stream_conv2d_4_source_20_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_20_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_20_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_20_pat_count_3 <= _source_stream_conv2d_4_source_20_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_20_source_pat_fsm_2 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_20_source_ram_renable <= 0;
        _stream_conv2d_4_source_20_idle <= 1;
      end 
      if((_stream_conv2d_4_source_20_source_pat_fsm_2 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_20_source_ram_renable <= 0;
        _stream_conv2d_4_source_20_idle <= 1;
      end 
      if(_set_flag_372) begin
        _stream_conv2d_4_source_21_source_mode <= 5'b10;
        _stream_conv2d_4_source_21_source_offset <= conv2d_4_stream_act_local_1 + conv2d_4_act_page_comp_offset_buf_0;
      end 
      if(_set_flag_372) begin
        _source_stream_conv2d_4_source_21_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_21_pat_stride_0 <= 1;
      end 
      if(_set_flag_372) begin
        _source_stream_conv2d_4_source_21_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_21_pat_stride_1 <= 0;
      end 
      if(_set_flag_372) begin
        _source_stream_conv2d_4_source_21_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_21_pat_stride_2 <= 0;
      end 
      if(_set_flag_372) begin
        _source_stream_conv2d_4_source_21_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_21_pat_stride_3 <= 0;
      end 
      if(_set_flag_372) begin
        _stream_conv2d_4_source_21_source_sel <= 4;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_21_source_offset_buf <= _stream_conv2d_4_source_21_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_count_0 <= _source_stream_conv2d_4_source_21_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_count_1 <= _source_stream_conv2d_4_source_21_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_count_2 <= _source_stream_conv2d_4_source_21_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_count_3 <= _source_stream_conv2d_4_source_21_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_size_buf_0 <= _source_stream_conv2d_4_source_21_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_size_buf_1 <= _source_stream_conv2d_4_source_21_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_size_buf_2 <= _source_stream_conv2d_4_source_21_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_size_buf_3 <= _source_stream_conv2d_4_source_21_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_stride_buf_0 <= _source_stream_conv2d_4_source_21_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_stride_buf_1 <= _source_stream_conv2d_4_source_21_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_stride_buf_2 <= _source_stream_conv2d_4_source_21_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_stride_buf_3 <= _source_stream_conv2d_4_source_21_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_1603 <= _stream_conv2d_4_source_21_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_21_source_pat_fsm_3 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_21_idle <= 0;
        _stream_conv2d_4_source_21_source_ram_raddr <= _stream_conv2d_4_source_21_source_pat_all_offset;
        _stream_conv2d_4_source_21_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_21_source_pat_fsm_3 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_cur_offset_0 <= _source_stream_conv2d_4_source_21_pat_cur_offset_0 + _source_stream_conv2d_4_source_21_pat_stride_buf_0;
        _source_stream_conv2d_4_source_21_pat_count_0 <= _source_stream_conv2d_4_source_21_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_21_source_pat_fsm_3 == 1) && (_source_stream_conv2d_4_source_21_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_21_pat_count_0 <= _source_stream_conv2d_4_source_21_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_21_source_pat_fsm_3 == 1) && (_source_stream_conv2d_4_source_21_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_cur_offset_1 <= _source_stream_conv2d_4_source_21_pat_cur_offset_1 + _source_stream_conv2d_4_source_21_pat_stride_buf_1;
        _source_stream_conv2d_4_source_21_pat_count_1 <= _source_stream_conv2d_4_source_21_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_21_source_pat_fsm_3 == 1) && (_source_stream_conv2d_4_source_21_pat_count_0 == 0) && (_source_stream_conv2d_4_source_21_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_21_pat_count_1 <= _source_stream_conv2d_4_source_21_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_21_source_pat_fsm_3 == 1) && ((_source_stream_conv2d_4_source_21_pat_count_0 == 0) && (_source_stream_conv2d_4_source_21_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_cur_offset_2 <= _source_stream_conv2d_4_source_21_pat_cur_offset_2 + _source_stream_conv2d_4_source_21_pat_stride_buf_2;
        _source_stream_conv2d_4_source_21_pat_count_2 <= _source_stream_conv2d_4_source_21_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_21_source_pat_fsm_3 == 1) && ((_source_stream_conv2d_4_source_21_pat_count_0 == 0) && (_source_stream_conv2d_4_source_21_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_21_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_21_pat_count_2 <= _source_stream_conv2d_4_source_21_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_21_source_pat_fsm_3 == 1) && ((_source_stream_conv2d_4_source_21_pat_count_0 == 0) && (_source_stream_conv2d_4_source_21_pat_count_1 == 0) && (_source_stream_conv2d_4_source_21_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_cur_offset_3 <= _source_stream_conv2d_4_source_21_pat_cur_offset_3 + _source_stream_conv2d_4_source_21_pat_stride_buf_3;
        _source_stream_conv2d_4_source_21_pat_count_3 <= _source_stream_conv2d_4_source_21_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_21_source_pat_fsm_3 == 1) && ((_source_stream_conv2d_4_source_21_pat_count_0 == 0) && (_source_stream_conv2d_4_source_21_pat_count_1 == 0) && (_source_stream_conv2d_4_source_21_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_21_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_21_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_21_pat_count_3 <= _source_stream_conv2d_4_source_21_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_21_source_pat_fsm_3 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_21_source_ram_renable <= 0;
        _stream_conv2d_4_source_21_idle <= 1;
      end 
      if((_stream_conv2d_4_source_21_source_pat_fsm_3 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_21_source_ram_renable <= 0;
        _stream_conv2d_4_source_21_idle <= 1;
      end 
      if(_set_flag_381) begin
        _stream_conv2d_4_source_22_source_mode <= 5'b10;
        _stream_conv2d_4_source_22_source_offset <= conv2d_4_stream_act_local_2 + conv2d_4_act_page_comp_offset_buf_0;
      end 
      if(_set_flag_381) begin
        _source_stream_conv2d_4_source_22_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_22_pat_stride_0 <= 1;
      end 
      if(_set_flag_381) begin
        _source_stream_conv2d_4_source_22_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_22_pat_stride_1 <= 0;
      end 
      if(_set_flag_381) begin
        _source_stream_conv2d_4_source_22_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_22_pat_stride_2 <= 0;
      end 
      if(_set_flag_381) begin
        _source_stream_conv2d_4_source_22_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_22_pat_stride_3 <= 0;
      end 
      if(_set_flag_381) begin
        _stream_conv2d_4_source_22_source_sel <= 5;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_22_source_offset_buf <= _stream_conv2d_4_source_22_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_count_0 <= _source_stream_conv2d_4_source_22_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_count_1 <= _source_stream_conv2d_4_source_22_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_count_2 <= _source_stream_conv2d_4_source_22_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_count_3 <= _source_stream_conv2d_4_source_22_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_size_buf_0 <= _source_stream_conv2d_4_source_22_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_size_buf_1 <= _source_stream_conv2d_4_source_22_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_size_buf_2 <= _source_stream_conv2d_4_source_22_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_size_buf_3 <= _source_stream_conv2d_4_source_22_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_stride_buf_0 <= _source_stream_conv2d_4_source_22_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_stride_buf_1 <= _source_stream_conv2d_4_source_22_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_stride_buf_2 <= _source_stream_conv2d_4_source_22_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_stride_buf_3 <= _source_stream_conv2d_4_source_22_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_1604 <= _stream_conv2d_4_source_22_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_22_source_pat_fsm_4 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_22_idle <= 0;
        _stream_conv2d_4_source_22_source_ram_raddr <= _stream_conv2d_4_source_22_source_pat_all_offset;
        _stream_conv2d_4_source_22_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_22_source_pat_fsm_4 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_cur_offset_0 <= _source_stream_conv2d_4_source_22_pat_cur_offset_0 + _source_stream_conv2d_4_source_22_pat_stride_buf_0;
        _source_stream_conv2d_4_source_22_pat_count_0 <= _source_stream_conv2d_4_source_22_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_22_source_pat_fsm_4 == 1) && (_source_stream_conv2d_4_source_22_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_22_pat_count_0 <= _source_stream_conv2d_4_source_22_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_22_source_pat_fsm_4 == 1) && (_source_stream_conv2d_4_source_22_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_cur_offset_1 <= _source_stream_conv2d_4_source_22_pat_cur_offset_1 + _source_stream_conv2d_4_source_22_pat_stride_buf_1;
        _source_stream_conv2d_4_source_22_pat_count_1 <= _source_stream_conv2d_4_source_22_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_22_source_pat_fsm_4 == 1) && (_source_stream_conv2d_4_source_22_pat_count_0 == 0) && (_source_stream_conv2d_4_source_22_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_22_pat_count_1 <= _source_stream_conv2d_4_source_22_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_22_source_pat_fsm_4 == 1) && ((_source_stream_conv2d_4_source_22_pat_count_0 == 0) && (_source_stream_conv2d_4_source_22_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_cur_offset_2 <= _source_stream_conv2d_4_source_22_pat_cur_offset_2 + _source_stream_conv2d_4_source_22_pat_stride_buf_2;
        _source_stream_conv2d_4_source_22_pat_count_2 <= _source_stream_conv2d_4_source_22_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_22_source_pat_fsm_4 == 1) && ((_source_stream_conv2d_4_source_22_pat_count_0 == 0) && (_source_stream_conv2d_4_source_22_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_22_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_22_pat_count_2 <= _source_stream_conv2d_4_source_22_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_22_source_pat_fsm_4 == 1) && ((_source_stream_conv2d_4_source_22_pat_count_0 == 0) && (_source_stream_conv2d_4_source_22_pat_count_1 == 0) && (_source_stream_conv2d_4_source_22_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_cur_offset_3 <= _source_stream_conv2d_4_source_22_pat_cur_offset_3 + _source_stream_conv2d_4_source_22_pat_stride_buf_3;
        _source_stream_conv2d_4_source_22_pat_count_3 <= _source_stream_conv2d_4_source_22_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_22_source_pat_fsm_4 == 1) && ((_source_stream_conv2d_4_source_22_pat_count_0 == 0) && (_source_stream_conv2d_4_source_22_pat_count_1 == 0) && (_source_stream_conv2d_4_source_22_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_22_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_22_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_22_pat_count_3 <= _source_stream_conv2d_4_source_22_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_22_source_pat_fsm_4 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_22_source_ram_renable <= 0;
        _stream_conv2d_4_source_22_idle <= 1;
      end 
      if((_stream_conv2d_4_source_22_source_pat_fsm_4 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_22_source_ram_renable <= 0;
        _stream_conv2d_4_source_22_idle <= 1;
      end 
      if(_set_flag_390) begin
        _stream_conv2d_4_source_23_source_mode <= 5'b10;
        _stream_conv2d_4_source_23_source_offset <= conv2d_4_stream_act_local_3 + conv2d_4_act_page_comp_offset_buf_1;
      end 
      if(_set_flag_390) begin
        _source_stream_conv2d_4_source_23_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_23_pat_stride_0 <= 1;
      end 
      if(_set_flag_390) begin
        _source_stream_conv2d_4_source_23_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_23_pat_stride_1 <= 0;
      end 
      if(_set_flag_390) begin
        _source_stream_conv2d_4_source_23_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_23_pat_stride_2 <= 0;
      end 
      if(_set_flag_390) begin
        _source_stream_conv2d_4_source_23_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_23_pat_stride_3 <= 0;
      end 
      if(_set_flag_390) begin
        _stream_conv2d_4_source_23_source_sel <= 6;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_23_source_offset_buf <= _stream_conv2d_4_source_23_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_count_0 <= _source_stream_conv2d_4_source_23_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_count_1 <= _source_stream_conv2d_4_source_23_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_count_2 <= _source_stream_conv2d_4_source_23_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_count_3 <= _source_stream_conv2d_4_source_23_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_size_buf_0 <= _source_stream_conv2d_4_source_23_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_size_buf_1 <= _source_stream_conv2d_4_source_23_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_size_buf_2 <= _source_stream_conv2d_4_source_23_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_size_buf_3 <= _source_stream_conv2d_4_source_23_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_stride_buf_0 <= _source_stream_conv2d_4_source_23_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_stride_buf_1 <= _source_stream_conv2d_4_source_23_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_stride_buf_2 <= _source_stream_conv2d_4_source_23_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_stride_buf_3 <= _source_stream_conv2d_4_source_23_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_1605 <= _stream_conv2d_4_source_23_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_23_source_pat_fsm_5 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_23_idle <= 0;
        _stream_conv2d_4_source_23_source_ram_raddr <= _stream_conv2d_4_source_23_source_pat_all_offset;
        _stream_conv2d_4_source_23_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_23_source_pat_fsm_5 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_cur_offset_0 <= _source_stream_conv2d_4_source_23_pat_cur_offset_0 + _source_stream_conv2d_4_source_23_pat_stride_buf_0;
        _source_stream_conv2d_4_source_23_pat_count_0 <= _source_stream_conv2d_4_source_23_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_23_source_pat_fsm_5 == 1) && (_source_stream_conv2d_4_source_23_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_23_pat_count_0 <= _source_stream_conv2d_4_source_23_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_23_source_pat_fsm_5 == 1) && (_source_stream_conv2d_4_source_23_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_cur_offset_1 <= _source_stream_conv2d_4_source_23_pat_cur_offset_1 + _source_stream_conv2d_4_source_23_pat_stride_buf_1;
        _source_stream_conv2d_4_source_23_pat_count_1 <= _source_stream_conv2d_4_source_23_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_23_source_pat_fsm_5 == 1) && (_source_stream_conv2d_4_source_23_pat_count_0 == 0) && (_source_stream_conv2d_4_source_23_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_23_pat_count_1 <= _source_stream_conv2d_4_source_23_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_23_source_pat_fsm_5 == 1) && ((_source_stream_conv2d_4_source_23_pat_count_0 == 0) && (_source_stream_conv2d_4_source_23_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_cur_offset_2 <= _source_stream_conv2d_4_source_23_pat_cur_offset_2 + _source_stream_conv2d_4_source_23_pat_stride_buf_2;
        _source_stream_conv2d_4_source_23_pat_count_2 <= _source_stream_conv2d_4_source_23_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_23_source_pat_fsm_5 == 1) && ((_source_stream_conv2d_4_source_23_pat_count_0 == 0) && (_source_stream_conv2d_4_source_23_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_23_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_23_pat_count_2 <= _source_stream_conv2d_4_source_23_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_23_source_pat_fsm_5 == 1) && ((_source_stream_conv2d_4_source_23_pat_count_0 == 0) && (_source_stream_conv2d_4_source_23_pat_count_1 == 0) && (_source_stream_conv2d_4_source_23_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_cur_offset_3 <= _source_stream_conv2d_4_source_23_pat_cur_offset_3 + _source_stream_conv2d_4_source_23_pat_stride_buf_3;
        _source_stream_conv2d_4_source_23_pat_count_3 <= _source_stream_conv2d_4_source_23_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_23_source_pat_fsm_5 == 1) && ((_source_stream_conv2d_4_source_23_pat_count_0 == 0) && (_source_stream_conv2d_4_source_23_pat_count_1 == 0) && (_source_stream_conv2d_4_source_23_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_23_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_23_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_23_pat_count_3 <= _source_stream_conv2d_4_source_23_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_23_source_pat_fsm_5 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_23_source_ram_renable <= 0;
        _stream_conv2d_4_source_23_idle <= 1;
      end 
      if((_stream_conv2d_4_source_23_source_pat_fsm_5 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_23_source_ram_renable <= 0;
        _stream_conv2d_4_source_23_idle <= 1;
      end 
      if(_set_flag_399) begin
        _stream_conv2d_4_source_24_source_mode <= 5'b10;
        _stream_conv2d_4_source_24_source_offset <= conv2d_4_stream_act_local_4 + conv2d_4_act_page_comp_offset_buf_1;
      end 
      if(_set_flag_399) begin
        _source_stream_conv2d_4_source_24_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_24_pat_stride_0 <= 1;
      end 
      if(_set_flag_399) begin
        _source_stream_conv2d_4_source_24_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_24_pat_stride_1 <= 0;
      end 
      if(_set_flag_399) begin
        _source_stream_conv2d_4_source_24_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_24_pat_stride_2 <= 0;
      end 
      if(_set_flag_399) begin
        _source_stream_conv2d_4_source_24_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_24_pat_stride_3 <= 0;
      end 
      if(_set_flag_399) begin
        _stream_conv2d_4_source_24_source_sel <= 7;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_24_source_offset_buf <= _stream_conv2d_4_source_24_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_count_0 <= _source_stream_conv2d_4_source_24_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_count_1 <= _source_stream_conv2d_4_source_24_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_count_2 <= _source_stream_conv2d_4_source_24_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_count_3 <= _source_stream_conv2d_4_source_24_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_size_buf_0 <= _source_stream_conv2d_4_source_24_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_size_buf_1 <= _source_stream_conv2d_4_source_24_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_size_buf_2 <= _source_stream_conv2d_4_source_24_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_size_buf_3 <= _source_stream_conv2d_4_source_24_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_stride_buf_0 <= _source_stream_conv2d_4_source_24_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_stride_buf_1 <= _source_stream_conv2d_4_source_24_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_stride_buf_2 <= _source_stream_conv2d_4_source_24_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_stride_buf_3 <= _source_stream_conv2d_4_source_24_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_1606 <= _stream_conv2d_4_source_24_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_24_source_pat_fsm_6 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_24_idle <= 0;
        _stream_conv2d_4_source_24_source_ram_raddr <= _stream_conv2d_4_source_24_source_pat_all_offset;
        _stream_conv2d_4_source_24_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_24_source_pat_fsm_6 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_cur_offset_0 <= _source_stream_conv2d_4_source_24_pat_cur_offset_0 + _source_stream_conv2d_4_source_24_pat_stride_buf_0;
        _source_stream_conv2d_4_source_24_pat_count_0 <= _source_stream_conv2d_4_source_24_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_24_source_pat_fsm_6 == 1) && (_source_stream_conv2d_4_source_24_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_24_pat_count_0 <= _source_stream_conv2d_4_source_24_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_24_source_pat_fsm_6 == 1) && (_source_stream_conv2d_4_source_24_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_cur_offset_1 <= _source_stream_conv2d_4_source_24_pat_cur_offset_1 + _source_stream_conv2d_4_source_24_pat_stride_buf_1;
        _source_stream_conv2d_4_source_24_pat_count_1 <= _source_stream_conv2d_4_source_24_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_24_source_pat_fsm_6 == 1) && (_source_stream_conv2d_4_source_24_pat_count_0 == 0) && (_source_stream_conv2d_4_source_24_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_24_pat_count_1 <= _source_stream_conv2d_4_source_24_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_24_source_pat_fsm_6 == 1) && ((_source_stream_conv2d_4_source_24_pat_count_0 == 0) && (_source_stream_conv2d_4_source_24_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_cur_offset_2 <= _source_stream_conv2d_4_source_24_pat_cur_offset_2 + _source_stream_conv2d_4_source_24_pat_stride_buf_2;
        _source_stream_conv2d_4_source_24_pat_count_2 <= _source_stream_conv2d_4_source_24_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_24_source_pat_fsm_6 == 1) && ((_source_stream_conv2d_4_source_24_pat_count_0 == 0) && (_source_stream_conv2d_4_source_24_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_24_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_24_pat_count_2 <= _source_stream_conv2d_4_source_24_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_24_source_pat_fsm_6 == 1) && ((_source_stream_conv2d_4_source_24_pat_count_0 == 0) && (_source_stream_conv2d_4_source_24_pat_count_1 == 0) && (_source_stream_conv2d_4_source_24_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_cur_offset_3 <= _source_stream_conv2d_4_source_24_pat_cur_offset_3 + _source_stream_conv2d_4_source_24_pat_stride_buf_3;
        _source_stream_conv2d_4_source_24_pat_count_3 <= _source_stream_conv2d_4_source_24_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_24_source_pat_fsm_6 == 1) && ((_source_stream_conv2d_4_source_24_pat_count_0 == 0) && (_source_stream_conv2d_4_source_24_pat_count_1 == 0) && (_source_stream_conv2d_4_source_24_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_24_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_24_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_24_pat_count_3 <= _source_stream_conv2d_4_source_24_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_24_source_pat_fsm_6 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_24_source_ram_renable <= 0;
        _stream_conv2d_4_source_24_idle <= 1;
      end 
      if((_stream_conv2d_4_source_24_source_pat_fsm_6 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_24_source_ram_renable <= 0;
        _stream_conv2d_4_source_24_idle <= 1;
      end 
      if(_set_flag_408) begin
        _stream_conv2d_4_source_25_source_mode <= 5'b10;
        _stream_conv2d_4_source_25_source_offset <= conv2d_4_stream_act_local_5 + conv2d_4_act_page_comp_offset_buf_1;
      end 
      if(_set_flag_408) begin
        _source_stream_conv2d_4_source_25_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_25_pat_stride_0 <= 1;
      end 
      if(_set_flag_408) begin
        _source_stream_conv2d_4_source_25_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_25_pat_stride_1 <= 0;
      end 
      if(_set_flag_408) begin
        _source_stream_conv2d_4_source_25_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_25_pat_stride_2 <= 0;
      end 
      if(_set_flag_408) begin
        _source_stream_conv2d_4_source_25_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_25_pat_stride_3 <= 0;
      end 
      if(_set_flag_408) begin
        _stream_conv2d_4_source_25_source_sel <= 8;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_25_source_offset_buf <= _stream_conv2d_4_source_25_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_count_0 <= _source_stream_conv2d_4_source_25_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_count_1 <= _source_stream_conv2d_4_source_25_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_count_2 <= _source_stream_conv2d_4_source_25_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_count_3 <= _source_stream_conv2d_4_source_25_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_size_buf_0 <= _source_stream_conv2d_4_source_25_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_size_buf_1 <= _source_stream_conv2d_4_source_25_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_size_buf_2 <= _source_stream_conv2d_4_source_25_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_size_buf_3 <= _source_stream_conv2d_4_source_25_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_stride_buf_0 <= _source_stream_conv2d_4_source_25_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_stride_buf_1 <= _source_stream_conv2d_4_source_25_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_stride_buf_2 <= _source_stream_conv2d_4_source_25_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_stride_buf_3 <= _source_stream_conv2d_4_source_25_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_1607 <= _stream_conv2d_4_source_25_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_25_source_pat_fsm_7 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_25_idle <= 0;
        _stream_conv2d_4_source_25_source_ram_raddr <= _stream_conv2d_4_source_25_source_pat_all_offset;
        _stream_conv2d_4_source_25_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_25_source_pat_fsm_7 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_cur_offset_0 <= _source_stream_conv2d_4_source_25_pat_cur_offset_0 + _source_stream_conv2d_4_source_25_pat_stride_buf_0;
        _source_stream_conv2d_4_source_25_pat_count_0 <= _source_stream_conv2d_4_source_25_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_25_source_pat_fsm_7 == 1) && (_source_stream_conv2d_4_source_25_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_25_pat_count_0 <= _source_stream_conv2d_4_source_25_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_25_source_pat_fsm_7 == 1) && (_source_stream_conv2d_4_source_25_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_cur_offset_1 <= _source_stream_conv2d_4_source_25_pat_cur_offset_1 + _source_stream_conv2d_4_source_25_pat_stride_buf_1;
        _source_stream_conv2d_4_source_25_pat_count_1 <= _source_stream_conv2d_4_source_25_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_25_source_pat_fsm_7 == 1) && (_source_stream_conv2d_4_source_25_pat_count_0 == 0) && (_source_stream_conv2d_4_source_25_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_25_pat_count_1 <= _source_stream_conv2d_4_source_25_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_25_source_pat_fsm_7 == 1) && ((_source_stream_conv2d_4_source_25_pat_count_0 == 0) && (_source_stream_conv2d_4_source_25_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_cur_offset_2 <= _source_stream_conv2d_4_source_25_pat_cur_offset_2 + _source_stream_conv2d_4_source_25_pat_stride_buf_2;
        _source_stream_conv2d_4_source_25_pat_count_2 <= _source_stream_conv2d_4_source_25_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_25_source_pat_fsm_7 == 1) && ((_source_stream_conv2d_4_source_25_pat_count_0 == 0) && (_source_stream_conv2d_4_source_25_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_25_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_25_pat_count_2 <= _source_stream_conv2d_4_source_25_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_25_source_pat_fsm_7 == 1) && ((_source_stream_conv2d_4_source_25_pat_count_0 == 0) && (_source_stream_conv2d_4_source_25_pat_count_1 == 0) && (_source_stream_conv2d_4_source_25_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_cur_offset_3 <= _source_stream_conv2d_4_source_25_pat_cur_offset_3 + _source_stream_conv2d_4_source_25_pat_stride_buf_3;
        _source_stream_conv2d_4_source_25_pat_count_3 <= _source_stream_conv2d_4_source_25_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_25_source_pat_fsm_7 == 1) && ((_source_stream_conv2d_4_source_25_pat_count_0 == 0) && (_source_stream_conv2d_4_source_25_pat_count_1 == 0) && (_source_stream_conv2d_4_source_25_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_25_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_25_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_25_pat_count_3 <= _source_stream_conv2d_4_source_25_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_25_source_pat_fsm_7 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_25_source_ram_renable <= 0;
        _stream_conv2d_4_source_25_idle <= 1;
      end 
      if((_stream_conv2d_4_source_25_source_pat_fsm_7 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_25_source_ram_renable <= 0;
        _stream_conv2d_4_source_25_idle <= 1;
      end 
      if(_set_flag_417) begin
        _stream_conv2d_4_source_26_source_mode <= 5'b10;
        _stream_conv2d_4_source_26_source_offset <= conv2d_4_stream_act_local_6 + conv2d_4_act_page_comp_offset_buf_2;
      end 
      if(_set_flag_417) begin
        _source_stream_conv2d_4_source_26_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_26_pat_stride_0 <= 1;
      end 
      if(_set_flag_417) begin
        _source_stream_conv2d_4_source_26_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_26_pat_stride_1 <= 0;
      end 
      if(_set_flag_417) begin
        _source_stream_conv2d_4_source_26_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_26_pat_stride_2 <= 0;
      end 
      if(_set_flag_417) begin
        _source_stream_conv2d_4_source_26_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_26_pat_stride_3 <= 0;
      end 
      if(_set_flag_417) begin
        _stream_conv2d_4_source_26_source_sel <= 9;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_26_source_offset_buf <= _stream_conv2d_4_source_26_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_count_0 <= _source_stream_conv2d_4_source_26_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_count_1 <= _source_stream_conv2d_4_source_26_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_count_2 <= _source_stream_conv2d_4_source_26_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_count_3 <= _source_stream_conv2d_4_source_26_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_size_buf_0 <= _source_stream_conv2d_4_source_26_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_size_buf_1 <= _source_stream_conv2d_4_source_26_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_size_buf_2 <= _source_stream_conv2d_4_source_26_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_size_buf_3 <= _source_stream_conv2d_4_source_26_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_stride_buf_0 <= _source_stream_conv2d_4_source_26_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_stride_buf_1 <= _source_stream_conv2d_4_source_26_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_stride_buf_2 <= _source_stream_conv2d_4_source_26_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_stride_buf_3 <= _source_stream_conv2d_4_source_26_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_1608 <= _stream_conv2d_4_source_26_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_26_source_pat_fsm_8 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_26_idle <= 0;
        _stream_conv2d_4_source_26_source_ram_raddr <= _stream_conv2d_4_source_26_source_pat_all_offset;
        _stream_conv2d_4_source_26_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_26_source_pat_fsm_8 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_cur_offset_0 <= _source_stream_conv2d_4_source_26_pat_cur_offset_0 + _source_stream_conv2d_4_source_26_pat_stride_buf_0;
        _source_stream_conv2d_4_source_26_pat_count_0 <= _source_stream_conv2d_4_source_26_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_26_source_pat_fsm_8 == 1) && (_source_stream_conv2d_4_source_26_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_26_pat_count_0 <= _source_stream_conv2d_4_source_26_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_26_source_pat_fsm_8 == 1) && (_source_stream_conv2d_4_source_26_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_cur_offset_1 <= _source_stream_conv2d_4_source_26_pat_cur_offset_1 + _source_stream_conv2d_4_source_26_pat_stride_buf_1;
        _source_stream_conv2d_4_source_26_pat_count_1 <= _source_stream_conv2d_4_source_26_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_26_source_pat_fsm_8 == 1) && (_source_stream_conv2d_4_source_26_pat_count_0 == 0) && (_source_stream_conv2d_4_source_26_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_26_pat_count_1 <= _source_stream_conv2d_4_source_26_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_26_source_pat_fsm_8 == 1) && ((_source_stream_conv2d_4_source_26_pat_count_0 == 0) && (_source_stream_conv2d_4_source_26_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_cur_offset_2 <= _source_stream_conv2d_4_source_26_pat_cur_offset_2 + _source_stream_conv2d_4_source_26_pat_stride_buf_2;
        _source_stream_conv2d_4_source_26_pat_count_2 <= _source_stream_conv2d_4_source_26_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_26_source_pat_fsm_8 == 1) && ((_source_stream_conv2d_4_source_26_pat_count_0 == 0) && (_source_stream_conv2d_4_source_26_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_26_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_26_pat_count_2 <= _source_stream_conv2d_4_source_26_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_26_source_pat_fsm_8 == 1) && ((_source_stream_conv2d_4_source_26_pat_count_0 == 0) && (_source_stream_conv2d_4_source_26_pat_count_1 == 0) && (_source_stream_conv2d_4_source_26_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_cur_offset_3 <= _source_stream_conv2d_4_source_26_pat_cur_offset_3 + _source_stream_conv2d_4_source_26_pat_stride_buf_3;
        _source_stream_conv2d_4_source_26_pat_count_3 <= _source_stream_conv2d_4_source_26_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_26_source_pat_fsm_8 == 1) && ((_source_stream_conv2d_4_source_26_pat_count_0 == 0) && (_source_stream_conv2d_4_source_26_pat_count_1 == 0) && (_source_stream_conv2d_4_source_26_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_26_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_26_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_26_pat_count_3 <= _source_stream_conv2d_4_source_26_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_26_source_pat_fsm_8 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_26_source_ram_renable <= 0;
        _stream_conv2d_4_source_26_idle <= 1;
      end 
      if((_stream_conv2d_4_source_26_source_pat_fsm_8 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_26_source_ram_renable <= 0;
        _stream_conv2d_4_source_26_idle <= 1;
      end 
      if(_set_flag_426) begin
        _stream_conv2d_4_source_27_source_mode <= 5'b10;
        _stream_conv2d_4_source_27_source_offset <= conv2d_4_stream_act_local_7 + conv2d_4_act_page_comp_offset_buf_2;
      end 
      if(_set_flag_426) begin
        _source_stream_conv2d_4_source_27_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_27_pat_stride_0 <= 1;
      end 
      if(_set_flag_426) begin
        _source_stream_conv2d_4_source_27_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_27_pat_stride_1 <= 0;
      end 
      if(_set_flag_426) begin
        _source_stream_conv2d_4_source_27_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_27_pat_stride_2 <= 0;
      end 
      if(_set_flag_426) begin
        _source_stream_conv2d_4_source_27_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_27_pat_stride_3 <= 0;
      end 
      if(_set_flag_426) begin
        _stream_conv2d_4_source_27_source_sel <= 10;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_27_source_offset_buf <= _stream_conv2d_4_source_27_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_count_0 <= _source_stream_conv2d_4_source_27_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_count_1 <= _source_stream_conv2d_4_source_27_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_count_2 <= _source_stream_conv2d_4_source_27_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_count_3 <= _source_stream_conv2d_4_source_27_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_size_buf_0 <= _source_stream_conv2d_4_source_27_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_size_buf_1 <= _source_stream_conv2d_4_source_27_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_size_buf_2 <= _source_stream_conv2d_4_source_27_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_size_buf_3 <= _source_stream_conv2d_4_source_27_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_stride_buf_0 <= _source_stream_conv2d_4_source_27_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_stride_buf_1 <= _source_stream_conv2d_4_source_27_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_stride_buf_2 <= _source_stream_conv2d_4_source_27_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_stride_buf_3 <= _source_stream_conv2d_4_source_27_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_1609 <= _stream_conv2d_4_source_27_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_27_source_pat_fsm_9 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_27_idle <= 0;
        _stream_conv2d_4_source_27_source_ram_raddr <= _stream_conv2d_4_source_27_source_pat_all_offset;
        _stream_conv2d_4_source_27_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_27_source_pat_fsm_9 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_cur_offset_0 <= _source_stream_conv2d_4_source_27_pat_cur_offset_0 + _source_stream_conv2d_4_source_27_pat_stride_buf_0;
        _source_stream_conv2d_4_source_27_pat_count_0 <= _source_stream_conv2d_4_source_27_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_27_source_pat_fsm_9 == 1) && (_source_stream_conv2d_4_source_27_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_27_pat_count_0 <= _source_stream_conv2d_4_source_27_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_27_source_pat_fsm_9 == 1) && (_source_stream_conv2d_4_source_27_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_cur_offset_1 <= _source_stream_conv2d_4_source_27_pat_cur_offset_1 + _source_stream_conv2d_4_source_27_pat_stride_buf_1;
        _source_stream_conv2d_4_source_27_pat_count_1 <= _source_stream_conv2d_4_source_27_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_27_source_pat_fsm_9 == 1) && (_source_stream_conv2d_4_source_27_pat_count_0 == 0) && (_source_stream_conv2d_4_source_27_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_27_pat_count_1 <= _source_stream_conv2d_4_source_27_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_27_source_pat_fsm_9 == 1) && ((_source_stream_conv2d_4_source_27_pat_count_0 == 0) && (_source_stream_conv2d_4_source_27_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_cur_offset_2 <= _source_stream_conv2d_4_source_27_pat_cur_offset_2 + _source_stream_conv2d_4_source_27_pat_stride_buf_2;
        _source_stream_conv2d_4_source_27_pat_count_2 <= _source_stream_conv2d_4_source_27_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_27_source_pat_fsm_9 == 1) && ((_source_stream_conv2d_4_source_27_pat_count_0 == 0) && (_source_stream_conv2d_4_source_27_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_27_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_27_pat_count_2 <= _source_stream_conv2d_4_source_27_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_27_source_pat_fsm_9 == 1) && ((_source_stream_conv2d_4_source_27_pat_count_0 == 0) && (_source_stream_conv2d_4_source_27_pat_count_1 == 0) && (_source_stream_conv2d_4_source_27_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_cur_offset_3 <= _source_stream_conv2d_4_source_27_pat_cur_offset_3 + _source_stream_conv2d_4_source_27_pat_stride_buf_3;
        _source_stream_conv2d_4_source_27_pat_count_3 <= _source_stream_conv2d_4_source_27_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_27_source_pat_fsm_9 == 1) && ((_source_stream_conv2d_4_source_27_pat_count_0 == 0) && (_source_stream_conv2d_4_source_27_pat_count_1 == 0) && (_source_stream_conv2d_4_source_27_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_27_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_27_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_27_pat_count_3 <= _source_stream_conv2d_4_source_27_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_27_source_pat_fsm_9 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_27_source_ram_renable <= 0;
        _stream_conv2d_4_source_27_idle <= 1;
      end 
      if((_stream_conv2d_4_source_27_source_pat_fsm_9 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_27_source_ram_renable <= 0;
        _stream_conv2d_4_source_27_idle <= 1;
      end 
      if(_set_flag_435) begin
        _stream_conv2d_4_source_28_source_mode <= 5'b10;
        _stream_conv2d_4_source_28_source_offset <= conv2d_4_stream_act_local_8 + conv2d_4_act_page_comp_offset_buf_2;
      end 
      if(_set_flag_435) begin
        _source_stream_conv2d_4_source_28_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_28_pat_stride_0 <= 1;
      end 
      if(_set_flag_435) begin
        _source_stream_conv2d_4_source_28_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_28_pat_stride_1 <= 0;
      end 
      if(_set_flag_435) begin
        _source_stream_conv2d_4_source_28_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_28_pat_stride_2 <= 0;
      end 
      if(_set_flag_435) begin
        _source_stream_conv2d_4_source_28_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_28_pat_stride_3 <= 0;
      end 
      if(_set_flag_435) begin
        _stream_conv2d_4_source_28_source_sel <= 11;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_28_source_offset_buf <= _stream_conv2d_4_source_28_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_count_0 <= _source_stream_conv2d_4_source_28_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_count_1 <= _source_stream_conv2d_4_source_28_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_count_2 <= _source_stream_conv2d_4_source_28_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_count_3 <= _source_stream_conv2d_4_source_28_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_size_buf_0 <= _source_stream_conv2d_4_source_28_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_size_buf_1 <= _source_stream_conv2d_4_source_28_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_size_buf_2 <= _source_stream_conv2d_4_source_28_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_size_buf_3 <= _source_stream_conv2d_4_source_28_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_stride_buf_0 <= _source_stream_conv2d_4_source_28_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_stride_buf_1 <= _source_stream_conv2d_4_source_28_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_stride_buf_2 <= _source_stream_conv2d_4_source_28_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_stride_buf_3 <= _source_stream_conv2d_4_source_28_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_1610 <= _stream_conv2d_4_source_28_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_28_source_pat_fsm_10 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_28_idle <= 0;
        _stream_conv2d_4_source_28_source_ram_raddr <= _stream_conv2d_4_source_28_source_pat_all_offset;
        _stream_conv2d_4_source_28_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_28_source_pat_fsm_10 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_cur_offset_0 <= _source_stream_conv2d_4_source_28_pat_cur_offset_0 + _source_stream_conv2d_4_source_28_pat_stride_buf_0;
        _source_stream_conv2d_4_source_28_pat_count_0 <= _source_stream_conv2d_4_source_28_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_28_source_pat_fsm_10 == 1) && (_source_stream_conv2d_4_source_28_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_28_pat_count_0 <= _source_stream_conv2d_4_source_28_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_28_source_pat_fsm_10 == 1) && (_source_stream_conv2d_4_source_28_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_cur_offset_1 <= _source_stream_conv2d_4_source_28_pat_cur_offset_1 + _source_stream_conv2d_4_source_28_pat_stride_buf_1;
        _source_stream_conv2d_4_source_28_pat_count_1 <= _source_stream_conv2d_4_source_28_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_28_source_pat_fsm_10 == 1) && (_source_stream_conv2d_4_source_28_pat_count_0 == 0) && (_source_stream_conv2d_4_source_28_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_28_pat_count_1 <= _source_stream_conv2d_4_source_28_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_28_source_pat_fsm_10 == 1) && ((_source_stream_conv2d_4_source_28_pat_count_0 == 0) && (_source_stream_conv2d_4_source_28_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_cur_offset_2 <= _source_stream_conv2d_4_source_28_pat_cur_offset_2 + _source_stream_conv2d_4_source_28_pat_stride_buf_2;
        _source_stream_conv2d_4_source_28_pat_count_2 <= _source_stream_conv2d_4_source_28_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_28_source_pat_fsm_10 == 1) && ((_source_stream_conv2d_4_source_28_pat_count_0 == 0) && (_source_stream_conv2d_4_source_28_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_28_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_28_pat_count_2 <= _source_stream_conv2d_4_source_28_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_28_source_pat_fsm_10 == 1) && ((_source_stream_conv2d_4_source_28_pat_count_0 == 0) && (_source_stream_conv2d_4_source_28_pat_count_1 == 0) && (_source_stream_conv2d_4_source_28_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_cur_offset_3 <= _source_stream_conv2d_4_source_28_pat_cur_offset_3 + _source_stream_conv2d_4_source_28_pat_stride_buf_3;
        _source_stream_conv2d_4_source_28_pat_count_3 <= _source_stream_conv2d_4_source_28_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_28_source_pat_fsm_10 == 1) && ((_source_stream_conv2d_4_source_28_pat_count_0 == 0) && (_source_stream_conv2d_4_source_28_pat_count_1 == 0) && (_source_stream_conv2d_4_source_28_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_28_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_28_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_28_pat_count_3 <= _source_stream_conv2d_4_source_28_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_28_source_pat_fsm_10 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_28_source_ram_renable <= 0;
        _stream_conv2d_4_source_28_idle <= 1;
      end 
      if((_stream_conv2d_4_source_28_source_pat_fsm_10 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_28_source_ram_renable <= 0;
        _stream_conv2d_4_source_28_idle <= 1;
      end 
      if(_set_flag_444) begin
        _stream_conv2d_4_source_29_source_mode <= 5'b10;
        _stream_conv2d_4_source_29_source_offset <= conv2d_4_filter_page_comp_offset_buf;
      end 
      if(_set_flag_444) begin
        _source_stream_conv2d_4_source_29_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_29_pat_stride_0 <= 1;
      end 
      if(_set_flag_444) begin
        _source_stream_conv2d_4_source_29_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_29_pat_stride_1 <= cparam_conv2d_4_stream_aligned_reduce_size;
      end 
      if(_set_flag_444) begin
        _source_stream_conv2d_4_source_29_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_29_pat_stride_2 <= 0;
      end 
      if(_set_flag_444) begin
        _source_stream_conv2d_4_source_29_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_29_pat_stride_3 <= 0;
      end 
      if(_set_flag_444) begin
        _stream_conv2d_4_source_29_source_sel <= 12;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_29_source_offset_buf <= _stream_conv2d_4_source_29_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_count_0 <= _source_stream_conv2d_4_source_29_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_count_1 <= _source_stream_conv2d_4_source_29_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_count_2 <= _source_stream_conv2d_4_source_29_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_count_3 <= _source_stream_conv2d_4_source_29_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_size_buf_0 <= _source_stream_conv2d_4_source_29_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_size_buf_1 <= _source_stream_conv2d_4_source_29_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_size_buf_2 <= _source_stream_conv2d_4_source_29_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_size_buf_3 <= _source_stream_conv2d_4_source_29_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_stride_buf_0 <= _source_stream_conv2d_4_source_29_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_stride_buf_1 <= _source_stream_conv2d_4_source_29_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_stride_buf_2 <= _source_stream_conv2d_4_source_29_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_stride_buf_3 <= _source_stream_conv2d_4_source_29_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_1836 <= _stream_conv2d_4_source_29_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_29_source_pat_fsm_11 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_29_idle <= 0;
        _stream_conv2d_4_source_29_source_ram_raddr <= _stream_conv2d_4_source_29_source_pat_all_offset;
        _stream_conv2d_4_source_29_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_29_source_pat_fsm_11 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_cur_offset_0 <= _source_stream_conv2d_4_source_29_pat_cur_offset_0 + _source_stream_conv2d_4_source_29_pat_stride_buf_0;
        _source_stream_conv2d_4_source_29_pat_count_0 <= _source_stream_conv2d_4_source_29_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_29_source_pat_fsm_11 == 1) && (_source_stream_conv2d_4_source_29_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_29_pat_count_0 <= _source_stream_conv2d_4_source_29_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_29_source_pat_fsm_11 == 1) && (_source_stream_conv2d_4_source_29_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_cur_offset_1 <= _source_stream_conv2d_4_source_29_pat_cur_offset_1 + _source_stream_conv2d_4_source_29_pat_stride_buf_1;
        _source_stream_conv2d_4_source_29_pat_count_1 <= _source_stream_conv2d_4_source_29_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_29_source_pat_fsm_11 == 1) && (_source_stream_conv2d_4_source_29_pat_count_0 == 0) && (_source_stream_conv2d_4_source_29_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_29_pat_count_1 <= _source_stream_conv2d_4_source_29_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_29_source_pat_fsm_11 == 1) && ((_source_stream_conv2d_4_source_29_pat_count_0 == 0) && (_source_stream_conv2d_4_source_29_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_cur_offset_2 <= _source_stream_conv2d_4_source_29_pat_cur_offset_2 + _source_stream_conv2d_4_source_29_pat_stride_buf_2;
        _source_stream_conv2d_4_source_29_pat_count_2 <= _source_stream_conv2d_4_source_29_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_29_source_pat_fsm_11 == 1) && ((_source_stream_conv2d_4_source_29_pat_count_0 == 0) && (_source_stream_conv2d_4_source_29_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_29_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_29_pat_count_2 <= _source_stream_conv2d_4_source_29_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_29_source_pat_fsm_11 == 1) && ((_source_stream_conv2d_4_source_29_pat_count_0 == 0) && (_source_stream_conv2d_4_source_29_pat_count_1 == 0) && (_source_stream_conv2d_4_source_29_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_cur_offset_3 <= _source_stream_conv2d_4_source_29_pat_cur_offset_3 + _source_stream_conv2d_4_source_29_pat_stride_buf_3;
        _source_stream_conv2d_4_source_29_pat_count_3 <= _source_stream_conv2d_4_source_29_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_29_source_pat_fsm_11 == 1) && ((_source_stream_conv2d_4_source_29_pat_count_0 == 0) && (_source_stream_conv2d_4_source_29_pat_count_1 == 0) && (_source_stream_conv2d_4_source_29_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_29_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_29_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_29_pat_count_3 <= _source_stream_conv2d_4_source_29_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_29_source_pat_fsm_11 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_29_source_ram_renable <= 0;
        _stream_conv2d_4_source_29_idle <= 1;
      end 
      if((_stream_conv2d_4_source_29_source_pat_fsm_11 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_29_source_ram_renable <= 0;
        _stream_conv2d_4_source_29_idle <= 1;
      end 
      if(_set_flag_453) begin
        _stream_conv2d_4_source_30_source_mode <= 5'b10;
        _stream_conv2d_4_source_30_source_offset <= conv2d_4_filter_page_comp_offset_buf;
      end 
      if(_set_flag_453) begin
        _source_stream_conv2d_4_source_30_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_30_pat_stride_0 <= 1;
      end 
      if(_set_flag_453) begin
        _source_stream_conv2d_4_source_30_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_30_pat_stride_1 <= cparam_conv2d_4_stream_aligned_reduce_size;
      end 
      if(_set_flag_453) begin
        _source_stream_conv2d_4_source_30_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_30_pat_stride_2 <= 0;
      end 
      if(_set_flag_453) begin
        _source_stream_conv2d_4_source_30_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_30_pat_stride_3 <= 0;
      end 
      if(_set_flag_453) begin
        _stream_conv2d_4_source_30_source_sel <= 13;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_30_source_offset_buf <= _stream_conv2d_4_source_30_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_count_0 <= _source_stream_conv2d_4_source_30_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_count_1 <= _source_stream_conv2d_4_source_30_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_count_2 <= _source_stream_conv2d_4_source_30_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_count_3 <= _source_stream_conv2d_4_source_30_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_size_buf_0 <= _source_stream_conv2d_4_source_30_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_size_buf_1 <= _source_stream_conv2d_4_source_30_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_size_buf_2 <= _source_stream_conv2d_4_source_30_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_size_buf_3 <= _source_stream_conv2d_4_source_30_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_stride_buf_0 <= _source_stream_conv2d_4_source_30_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_stride_buf_1 <= _source_stream_conv2d_4_source_30_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_stride_buf_2 <= _source_stream_conv2d_4_source_30_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_stride_buf_3 <= _source_stream_conv2d_4_source_30_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_1837 <= _stream_conv2d_4_source_30_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_30_source_pat_fsm_12 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_30_idle <= 0;
        _stream_conv2d_4_source_30_source_ram_raddr <= _stream_conv2d_4_source_30_source_pat_all_offset;
        _stream_conv2d_4_source_30_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_30_source_pat_fsm_12 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_cur_offset_0 <= _source_stream_conv2d_4_source_30_pat_cur_offset_0 + _source_stream_conv2d_4_source_30_pat_stride_buf_0;
        _source_stream_conv2d_4_source_30_pat_count_0 <= _source_stream_conv2d_4_source_30_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_30_source_pat_fsm_12 == 1) && (_source_stream_conv2d_4_source_30_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_30_pat_count_0 <= _source_stream_conv2d_4_source_30_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_30_source_pat_fsm_12 == 1) && (_source_stream_conv2d_4_source_30_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_cur_offset_1 <= _source_stream_conv2d_4_source_30_pat_cur_offset_1 + _source_stream_conv2d_4_source_30_pat_stride_buf_1;
        _source_stream_conv2d_4_source_30_pat_count_1 <= _source_stream_conv2d_4_source_30_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_30_source_pat_fsm_12 == 1) && (_source_stream_conv2d_4_source_30_pat_count_0 == 0) && (_source_stream_conv2d_4_source_30_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_30_pat_count_1 <= _source_stream_conv2d_4_source_30_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_30_source_pat_fsm_12 == 1) && ((_source_stream_conv2d_4_source_30_pat_count_0 == 0) && (_source_stream_conv2d_4_source_30_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_cur_offset_2 <= _source_stream_conv2d_4_source_30_pat_cur_offset_2 + _source_stream_conv2d_4_source_30_pat_stride_buf_2;
        _source_stream_conv2d_4_source_30_pat_count_2 <= _source_stream_conv2d_4_source_30_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_30_source_pat_fsm_12 == 1) && ((_source_stream_conv2d_4_source_30_pat_count_0 == 0) && (_source_stream_conv2d_4_source_30_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_30_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_30_pat_count_2 <= _source_stream_conv2d_4_source_30_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_30_source_pat_fsm_12 == 1) && ((_source_stream_conv2d_4_source_30_pat_count_0 == 0) && (_source_stream_conv2d_4_source_30_pat_count_1 == 0) && (_source_stream_conv2d_4_source_30_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_cur_offset_3 <= _source_stream_conv2d_4_source_30_pat_cur_offset_3 + _source_stream_conv2d_4_source_30_pat_stride_buf_3;
        _source_stream_conv2d_4_source_30_pat_count_3 <= _source_stream_conv2d_4_source_30_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_30_source_pat_fsm_12 == 1) && ((_source_stream_conv2d_4_source_30_pat_count_0 == 0) && (_source_stream_conv2d_4_source_30_pat_count_1 == 0) && (_source_stream_conv2d_4_source_30_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_30_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_30_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_30_pat_count_3 <= _source_stream_conv2d_4_source_30_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_30_source_pat_fsm_12 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_30_source_ram_renable <= 0;
        _stream_conv2d_4_source_30_idle <= 1;
      end 
      if((_stream_conv2d_4_source_30_source_pat_fsm_12 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_30_source_ram_renable <= 0;
        _stream_conv2d_4_source_30_idle <= 1;
      end 
      if(_set_flag_462) begin
        _stream_conv2d_4_source_31_source_mode <= 5'b10;
        _stream_conv2d_4_source_31_source_offset <= conv2d_4_filter_page_comp_offset_buf;
      end 
      if(_set_flag_462) begin
        _source_stream_conv2d_4_source_31_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_31_pat_stride_0 <= 1;
      end 
      if(_set_flag_462) begin
        _source_stream_conv2d_4_source_31_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_31_pat_stride_1 <= cparam_conv2d_4_stream_aligned_reduce_size;
      end 
      if(_set_flag_462) begin
        _source_stream_conv2d_4_source_31_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_31_pat_stride_2 <= 0;
      end 
      if(_set_flag_462) begin
        _source_stream_conv2d_4_source_31_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_31_pat_stride_3 <= 0;
      end 
      if(_set_flag_462) begin
        _stream_conv2d_4_source_31_source_sel <= 14;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_31_source_offset_buf <= _stream_conv2d_4_source_31_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_count_0 <= _source_stream_conv2d_4_source_31_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_count_1 <= _source_stream_conv2d_4_source_31_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_count_2 <= _source_stream_conv2d_4_source_31_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_count_3 <= _source_stream_conv2d_4_source_31_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_size_buf_0 <= _source_stream_conv2d_4_source_31_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_size_buf_1 <= _source_stream_conv2d_4_source_31_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_size_buf_2 <= _source_stream_conv2d_4_source_31_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_size_buf_3 <= _source_stream_conv2d_4_source_31_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_stride_buf_0 <= _source_stream_conv2d_4_source_31_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_stride_buf_1 <= _source_stream_conv2d_4_source_31_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_stride_buf_2 <= _source_stream_conv2d_4_source_31_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_stride_buf_3 <= _source_stream_conv2d_4_source_31_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_1838 <= _stream_conv2d_4_source_31_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_31_source_pat_fsm_13 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_31_idle <= 0;
        _stream_conv2d_4_source_31_source_ram_raddr <= _stream_conv2d_4_source_31_source_pat_all_offset;
        _stream_conv2d_4_source_31_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_31_source_pat_fsm_13 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_cur_offset_0 <= _source_stream_conv2d_4_source_31_pat_cur_offset_0 + _source_stream_conv2d_4_source_31_pat_stride_buf_0;
        _source_stream_conv2d_4_source_31_pat_count_0 <= _source_stream_conv2d_4_source_31_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_31_source_pat_fsm_13 == 1) && (_source_stream_conv2d_4_source_31_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_31_pat_count_0 <= _source_stream_conv2d_4_source_31_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_31_source_pat_fsm_13 == 1) && (_source_stream_conv2d_4_source_31_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_cur_offset_1 <= _source_stream_conv2d_4_source_31_pat_cur_offset_1 + _source_stream_conv2d_4_source_31_pat_stride_buf_1;
        _source_stream_conv2d_4_source_31_pat_count_1 <= _source_stream_conv2d_4_source_31_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_31_source_pat_fsm_13 == 1) && (_source_stream_conv2d_4_source_31_pat_count_0 == 0) && (_source_stream_conv2d_4_source_31_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_31_pat_count_1 <= _source_stream_conv2d_4_source_31_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_31_source_pat_fsm_13 == 1) && ((_source_stream_conv2d_4_source_31_pat_count_0 == 0) && (_source_stream_conv2d_4_source_31_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_cur_offset_2 <= _source_stream_conv2d_4_source_31_pat_cur_offset_2 + _source_stream_conv2d_4_source_31_pat_stride_buf_2;
        _source_stream_conv2d_4_source_31_pat_count_2 <= _source_stream_conv2d_4_source_31_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_31_source_pat_fsm_13 == 1) && ((_source_stream_conv2d_4_source_31_pat_count_0 == 0) && (_source_stream_conv2d_4_source_31_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_31_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_31_pat_count_2 <= _source_stream_conv2d_4_source_31_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_31_source_pat_fsm_13 == 1) && ((_source_stream_conv2d_4_source_31_pat_count_0 == 0) && (_source_stream_conv2d_4_source_31_pat_count_1 == 0) && (_source_stream_conv2d_4_source_31_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_cur_offset_3 <= _source_stream_conv2d_4_source_31_pat_cur_offset_3 + _source_stream_conv2d_4_source_31_pat_stride_buf_3;
        _source_stream_conv2d_4_source_31_pat_count_3 <= _source_stream_conv2d_4_source_31_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_31_source_pat_fsm_13 == 1) && ((_source_stream_conv2d_4_source_31_pat_count_0 == 0) && (_source_stream_conv2d_4_source_31_pat_count_1 == 0) && (_source_stream_conv2d_4_source_31_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_31_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_31_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_31_pat_count_3 <= _source_stream_conv2d_4_source_31_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_31_source_pat_fsm_13 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_31_source_ram_renable <= 0;
        _stream_conv2d_4_source_31_idle <= 1;
      end 
      if((_stream_conv2d_4_source_31_source_pat_fsm_13 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_31_source_ram_renable <= 0;
        _stream_conv2d_4_source_31_idle <= 1;
      end 
      if(_set_flag_471) begin
        _stream_conv2d_4_source_32_source_mode <= 5'b10;
        _stream_conv2d_4_source_32_source_offset <= conv2d_4_filter_page_comp_offset_buf;
      end 
      if(_set_flag_471) begin
        _source_stream_conv2d_4_source_32_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_32_pat_stride_0 <= 1;
      end 
      if(_set_flag_471) begin
        _source_stream_conv2d_4_source_32_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_32_pat_stride_1 <= cparam_conv2d_4_stream_aligned_reduce_size;
      end 
      if(_set_flag_471) begin
        _source_stream_conv2d_4_source_32_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_32_pat_stride_2 <= 0;
      end 
      if(_set_flag_471) begin
        _source_stream_conv2d_4_source_32_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_32_pat_stride_3 <= 0;
      end 
      if(_set_flag_471) begin
        _stream_conv2d_4_source_32_source_sel <= 15;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_32_source_offset_buf <= _stream_conv2d_4_source_32_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_count_0 <= _source_stream_conv2d_4_source_32_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_count_1 <= _source_stream_conv2d_4_source_32_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_count_2 <= _source_stream_conv2d_4_source_32_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_count_3 <= _source_stream_conv2d_4_source_32_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_size_buf_0 <= _source_stream_conv2d_4_source_32_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_size_buf_1 <= _source_stream_conv2d_4_source_32_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_size_buf_2 <= _source_stream_conv2d_4_source_32_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_size_buf_3 <= _source_stream_conv2d_4_source_32_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_stride_buf_0 <= _source_stream_conv2d_4_source_32_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_stride_buf_1 <= _source_stream_conv2d_4_source_32_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_stride_buf_2 <= _source_stream_conv2d_4_source_32_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_stride_buf_3 <= _source_stream_conv2d_4_source_32_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_1839 <= _stream_conv2d_4_source_32_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_32_source_pat_fsm_14 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_32_idle <= 0;
        _stream_conv2d_4_source_32_source_ram_raddr <= _stream_conv2d_4_source_32_source_pat_all_offset;
        _stream_conv2d_4_source_32_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_32_source_pat_fsm_14 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_cur_offset_0 <= _source_stream_conv2d_4_source_32_pat_cur_offset_0 + _source_stream_conv2d_4_source_32_pat_stride_buf_0;
        _source_stream_conv2d_4_source_32_pat_count_0 <= _source_stream_conv2d_4_source_32_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_32_source_pat_fsm_14 == 1) && (_source_stream_conv2d_4_source_32_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_32_pat_count_0 <= _source_stream_conv2d_4_source_32_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_32_source_pat_fsm_14 == 1) && (_source_stream_conv2d_4_source_32_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_cur_offset_1 <= _source_stream_conv2d_4_source_32_pat_cur_offset_1 + _source_stream_conv2d_4_source_32_pat_stride_buf_1;
        _source_stream_conv2d_4_source_32_pat_count_1 <= _source_stream_conv2d_4_source_32_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_32_source_pat_fsm_14 == 1) && (_source_stream_conv2d_4_source_32_pat_count_0 == 0) && (_source_stream_conv2d_4_source_32_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_32_pat_count_1 <= _source_stream_conv2d_4_source_32_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_32_source_pat_fsm_14 == 1) && ((_source_stream_conv2d_4_source_32_pat_count_0 == 0) && (_source_stream_conv2d_4_source_32_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_cur_offset_2 <= _source_stream_conv2d_4_source_32_pat_cur_offset_2 + _source_stream_conv2d_4_source_32_pat_stride_buf_2;
        _source_stream_conv2d_4_source_32_pat_count_2 <= _source_stream_conv2d_4_source_32_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_32_source_pat_fsm_14 == 1) && ((_source_stream_conv2d_4_source_32_pat_count_0 == 0) && (_source_stream_conv2d_4_source_32_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_32_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_32_pat_count_2 <= _source_stream_conv2d_4_source_32_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_32_source_pat_fsm_14 == 1) && ((_source_stream_conv2d_4_source_32_pat_count_0 == 0) && (_source_stream_conv2d_4_source_32_pat_count_1 == 0) && (_source_stream_conv2d_4_source_32_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_cur_offset_3 <= _source_stream_conv2d_4_source_32_pat_cur_offset_3 + _source_stream_conv2d_4_source_32_pat_stride_buf_3;
        _source_stream_conv2d_4_source_32_pat_count_3 <= _source_stream_conv2d_4_source_32_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_32_source_pat_fsm_14 == 1) && ((_source_stream_conv2d_4_source_32_pat_count_0 == 0) && (_source_stream_conv2d_4_source_32_pat_count_1 == 0) && (_source_stream_conv2d_4_source_32_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_32_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_32_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_32_pat_count_3 <= _source_stream_conv2d_4_source_32_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_32_source_pat_fsm_14 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_32_source_ram_renable <= 0;
        _stream_conv2d_4_source_32_idle <= 1;
      end 
      if((_stream_conv2d_4_source_32_source_pat_fsm_14 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_32_source_ram_renable <= 0;
        _stream_conv2d_4_source_32_idle <= 1;
      end 
      if(_set_flag_480) begin
        _stream_conv2d_4_source_33_source_mode <= 5'b10;
        _stream_conv2d_4_source_33_source_offset <= conv2d_4_filter_page_comp_offset_buf;
      end 
      if(_set_flag_480) begin
        _source_stream_conv2d_4_source_33_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_33_pat_stride_0 <= 1;
      end 
      if(_set_flag_480) begin
        _source_stream_conv2d_4_source_33_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_33_pat_stride_1 <= cparam_conv2d_4_stream_aligned_reduce_size;
      end 
      if(_set_flag_480) begin
        _source_stream_conv2d_4_source_33_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_33_pat_stride_2 <= 0;
      end 
      if(_set_flag_480) begin
        _source_stream_conv2d_4_source_33_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_33_pat_stride_3 <= 0;
      end 
      if(_set_flag_480) begin
        _stream_conv2d_4_source_33_source_sel <= 16;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_33_source_offset_buf <= _stream_conv2d_4_source_33_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_count_0 <= _source_stream_conv2d_4_source_33_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_count_1 <= _source_stream_conv2d_4_source_33_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_count_2 <= _source_stream_conv2d_4_source_33_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_count_3 <= _source_stream_conv2d_4_source_33_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_size_buf_0 <= _source_stream_conv2d_4_source_33_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_size_buf_1 <= _source_stream_conv2d_4_source_33_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_size_buf_2 <= _source_stream_conv2d_4_source_33_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_size_buf_3 <= _source_stream_conv2d_4_source_33_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_stride_buf_0 <= _source_stream_conv2d_4_source_33_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_stride_buf_1 <= _source_stream_conv2d_4_source_33_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_stride_buf_2 <= _source_stream_conv2d_4_source_33_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_stride_buf_3 <= _source_stream_conv2d_4_source_33_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_1840 <= _stream_conv2d_4_source_33_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_33_source_pat_fsm_15 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_33_idle <= 0;
        _stream_conv2d_4_source_33_source_ram_raddr <= _stream_conv2d_4_source_33_source_pat_all_offset;
        _stream_conv2d_4_source_33_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_33_source_pat_fsm_15 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_cur_offset_0 <= _source_stream_conv2d_4_source_33_pat_cur_offset_0 + _source_stream_conv2d_4_source_33_pat_stride_buf_0;
        _source_stream_conv2d_4_source_33_pat_count_0 <= _source_stream_conv2d_4_source_33_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_33_source_pat_fsm_15 == 1) && (_source_stream_conv2d_4_source_33_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_33_pat_count_0 <= _source_stream_conv2d_4_source_33_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_33_source_pat_fsm_15 == 1) && (_source_stream_conv2d_4_source_33_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_cur_offset_1 <= _source_stream_conv2d_4_source_33_pat_cur_offset_1 + _source_stream_conv2d_4_source_33_pat_stride_buf_1;
        _source_stream_conv2d_4_source_33_pat_count_1 <= _source_stream_conv2d_4_source_33_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_33_source_pat_fsm_15 == 1) && (_source_stream_conv2d_4_source_33_pat_count_0 == 0) && (_source_stream_conv2d_4_source_33_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_33_pat_count_1 <= _source_stream_conv2d_4_source_33_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_33_source_pat_fsm_15 == 1) && ((_source_stream_conv2d_4_source_33_pat_count_0 == 0) && (_source_stream_conv2d_4_source_33_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_cur_offset_2 <= _source_stream_conv2d_4_source_33_pat_cur_offset_2 + _source_stream_conv2d_4_source_33_pat_stride_buf_2;
        _source_stream_conv2d_4_source_33_pat_count_2 <= _source_stream_conv2d_4_source_33_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_33_source_pat_fsm_15 == 1) && ((_source_stream_conv2d_4_source_33_pat_count_0 == 0) && (_source_stream_conv2d_4_source_33_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_33_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_33_pat_count_2 <= _source_stream_conv2d_4_source_33_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_33_source_pat_fsm_15 == 1) && ((_source_stream_conv2d_4_source_33_pat_count_0 == 0) && (_source_stream_conv2d_4_source_33_pat_count_1 == 0) && (_source_stream_conv2d_4_source_33_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_cur_offset_3 <= _source_stream_conv2d_4_source_33_pat_cur_offset_3 + _source_stream_conv2d_4_source_33_pat_stride_buf_3;
        _source_stream_conv2d_4_source_33_pat_count_3 <= _source_stream_conv2d_4_source_33_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_33_source_pat_fsm_15 == 1) && ((_source_stream_conv2d_4_source_33_pat_count_0 == 0) && (_source_stream_conv2d_4_source_33_pat_count_1 == 0) && (_source_stream_conv2d_4_source_33_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_33_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_33_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_33_pat_count_3 <= _source_stream_conv2d_4_source_33_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_33_source_pat_fsm_15 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_33_source_ram_renable <= 0;
        _stream_conv2d_4_source_33_idle <= 1;
      end 
      if((_stream_conv2d_4_source_33_source_pat_fsm_15 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_33_source_ram_renable <= 0;
        _stream_conv2d_4_source_33_idle <= 1;
      end 
      if(_set_flag_489) begin
        _stream_conv2d_4_source_34_source_mode <= 5'b10;
        _stream_conv2d_4_source_34_source_offset <= conv2d_4_filter_page_comp_offset_buf;
      end 
      if(_set_flag_489) begin
        _source_stream_conv2d_4_source_34_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_34_pat_stride_0 <= 1;
      end 
      if(_set_flag_489) begin
        _source_stream_conv2d_4_source_34_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_34_pat_stride_1 <= cparam_conv2d_4_stream_aligned_reduce_size;
      end 
      if(_set_flag_489) begin
        _source_stream_conv2d_4_source_34_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_34_pat_stride_2 <= 0;
      end 
      if(_set_flag_489) begin
        _source_stream_conv2d_4_source_34_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_34_pat_stride_3 <= 0;
      end 
      if(_set_flag_489) begin
        _stream_conv2d_4_source_34_source_sel <= 17;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_34_source_offset_buf <= _stream_conv2d_4_source_34_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_count_0 <= _source_stream_conv2d_4_source_34_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_count_1 <= _source_stream_conv2d_4_source_34_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_count_2 <= _source_stream_conv2d_4_source_34_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_count_3 <= _source_stream_conv2d_4_source_34_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_size_buf_0 <= _source_stream_conv2d_4_source_34_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_size_buf_1 <= _source_stream_conv2d_4_source_34_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_size_buf_2 <= _source_stream_conv2d_4_source_34_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_size_buf_3 <= _source_stream_conv2d_4_source_34_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_stride_buf_0 <= _source_stream_conv2d_4_source_34_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_stride_buf_1 <= _source_stream_conv2d_4_source_34_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_stride_buf_2 <= _source_stream_conv2d_4_source_34_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_stride_buf_3 <= _source_stream_conv2d_4_source_34_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_1841 <= _stream_conv2d_4_source_34_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_34_source_pat_fsm_16 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_34_idle <= 0;
        _stream_conv2d_4_source_34_source_ram_raddr <= _stream_conv2d_4_source_34_source_pat_all_offset;
        _stream_conv2d_4_source_34_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_34_source_pat_fsm_16 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_cur_offset_0 <= _source_stream_conv2d_4_source_34_pat_cur_offset_0 + _source_stream_conv2d_4_source_34_pat_stride_buf_0;
        _source_stream_conv2d_4_source_34_pat_count_0 <= _source_stream_conv2d_4_source_34_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_34_source_pat_fsm_16 == 1) && (_source_stream_conv2d_4_source_34_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_34_pat_count_0 <= _source_stream_conv2d_4_source_34_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_34_source_pat_fsm_16 == 1) && (_source_stream_conv2d_4_source_34_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_cur_offset_1 <= _source_stream_conv2d_4_source_34_pat_cur_offset_1 + _source_stream_conv2d_4_source_34_pat_stride_buf_1;
        _source_stream_conv2d_4_source_34_pat_count_1 <= _source_stream_conv2d_4_source_34_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_34_source_pat_fsm_16 == 1) && (_source_stream_conv2d_4_source_34_pat_count_0 == 0) && (_source_stream_conv2d_4_source_34_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_34_pat_count_1 <= _source_stream_conv2d_4_source_34_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_34_source_pat_fsm_16 == 1) && ((_source_stream_conv2d_4_source_34_pat_count_0 == 0) && (_source_stream_conv2d_4_source_34_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_cur_offset_2 <= _source_stream_conv2d_4_source_34_pat_cur_offset_2 + _source_stream_conv2d_4_source_34_pat_stride_buf_2;
        _source_stream_conv2d_4_source_34_pat_count_2 <= _source_stream_conv2d_4_source_34_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_34_source_pat_fsm_16 == 1) && ((_source_stream_conv2d_4_source_34_pat_count_0 == 0) && (_source_stream_conv2d_4_source_34_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_34_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_34_pat_count_2 <= _source_stream_conv2d_4_source_34_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_34_source_pat_fsm_16 == 1) && ((_source_stream_conv2d_4_source_34_pat_count_0 == 0) && (_source_stream_conv2d_4_source_34_pat_count_1 == 0) && (_source_stream_conv2d_4_source_34_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_cur_offset_3 <= _source_stream_conv2d_4_source_34_pat_cur_offset_3 + _source_stream_conv2d_4_source_34_pat_stride_buf_3;
        _source_stream_conv2d_4_source_34_pat_count_3 <= _source_stream_conv2d_4_source_34_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_34_source_pat_fsm_16 == 1) && ((_source_stream_conv2d_4_source_34_pat_count_0 == 0) && (_source_stream_conv2d_4_source_34_pat_count_1 == 0) && (_source_stream_conv2d_4_source_34_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_34_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_34_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_34_pat_count_3 <= _source_stream_conv2d_4_source_34_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_34_source_pat_fsm_16 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_34_source_ram_renable <= 0;
        _stream_conv2d_4_source_34_idle <= 1;
      end 
      if((_stream_conv2d_4_source_34_source_pat_fsm_16 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_34_source_ram_renable <= 0;
        _stream_conv2d_4_source_34_idle <= 1;
      end 
      if(_set_flag_498) begin
        _stream_conv2d_4_source_35_source_mode <= 5'b10;
        _stream_conv2d_4_source_35_source_offset <= conv2d_4_filter_page_comp_offset_buf;
      end 
      if(_set_flag_498) begin
        _source_stream_conv2d_4_source_35_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_35_pat_stride_0 <= 1;
      end 
      if(_set_flag_498) begin
        _source_stream_conv2d_4_source_35_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_35_pat_stride_1 <= cparam_conv2d_4_stream_aligned_reduce_size;
      end 
      if(_set_flag_498) begin
        _source_stream_conv2d_4_source_35_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_35_pat_stride_2 <= 0;
      end 
      if(_set_flag_498) begin
        _source_stream_conv2d_4_source_35_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_35_pat_stride_3 <= 0;
      end 
      if(_set_flag_498) begin
        _stream_conv2d_4_source_35_source_sel <= 18;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_35_source_offset_buf <= _stream_conv2d_4_source_35_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_count_0 <= _source_stream_conv2d_4_source_35_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_count_1 <= _source_stream_conv2d_4_source_35_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_count_2 <= _source_stream_conv2d_4_source_35_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_count_3 <= _source_stream_conv2d_4_source_35_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_size_buf_0 <= _source_stream_conv2d_4_source_35_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_size_buf_1 <= _source_stream_conv2d_4_source_35_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_size_buf_2 <= _source_stream_conv2d_4_source_35_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_size_buf_3 <= _source_stream_conv2d_4_source_35_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_stride_buf_0 <= _source_stream_conv2d_4_source_35_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_stride_buf_1 <= _source_stream_conv2d_4_source_35_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_stride_buf_2 <= _source_stream_conv2d_4_source_35_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_stride_buf_3 <= _source_stream_conv2d_4_source_35_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_1842 <= _stream_conv2d_4_source_35_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_35_source_pat_fsm_17 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_35_idle <= 0;
        _stream_conv2d_4_source_35_source_ram_raddr <= _stream_conv2d_4_source_35_source_pat_all_offset;
        _stream_conv2d_4_source_35_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_35_source_pat_fsm_17 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_cur_offset_0 <= _source_stream_conv2d_4_source_35_pat_cur_offset_0 + _source_stream_conv2d_4_source_35_pat_stride_buf_0;
        _source_stream_conv2d_4_source_35_pat_count_0 <= _source_stream_conv2d_4_source_35_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_35_source_pat_fsm_17 == 1) && (_source_stream_conv2d_4_source_35_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_35_pat_count_0 <= _source_stream_conv2d_4_source_35_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_35_source_pat_fsm_17 == 1) && (_source_stream_conv2d_4_source_35_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_cur_offset_1 <= _source_stream_conv2d_4_source_35_pat_cur_offset_1 + _source_stream_conv2d_4_source_35_pat_stride_buf_1;
        _source_stream_conv2d_4_source_35_pat_count_1 <= _source_stream_conv2d_4_source_35_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_35_source_pat_fsm_17 == 1) && (_source_stream_conv2d_4_source_35_pat_count_0 == 0) && (_source_stream_conv2d_4_source_35_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_35_pat_count_1 <= _source_stream_conv2d_4_source_35_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_35_source_pat_fsm_17 == 1) && ((_source_stream_conv2d_4_source_35_pat_count_0 == 0) && (_source_stream_conv2d_4_source_35_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_cur_offset_2 <= _source_stream_conv2d_4_source_35_pat_cur_offset_2 + _source_stream_conv2d_4_source_35_pat_stride_buf_2;
        _source_stream_conv2d_4_source_35_pat_count_2 <= _source_stream_conv2d_4_source_35_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_35_source_pat_fsm_17 == 1) && ((_source_stream_conv2d_4_source_35_pat_count_0 == 0) && (_source_stream_conv2d_4_source_35_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_35_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_35_pat_count_2 <= _source_stream_conv2d_4_source_35_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_35_source_pat_fsm_17 == 1) && ((_source_stream_conv2d_4_source_35_pat_count_0 == 0) && (_source_stream_conv2d_4_source_35_pat_count_1 == 0) && (_source_stream_conv2d_4_source_35_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_cur_offset_3 <= _source_stream_conv2d_4_source_35_pat_cur_offset_3 + _source_stream_conv2d_4_source_35_pat_stride_buf_3;
        _source_stream_conv2d_4_source_35_pat_count_3 <= _source_stream_conv2d_4_source_35_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_35_source_pat_fsm_17 == 1) && ((_source_stream_conv2d_4_source_35_pat_count_0 == 0) && (_source_stream_conv2d_4_source_35_pat_count_1 == 0) && (_source_stream_conv2d_4_source_35_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_35_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_35_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_35_pat_count_3 <= _source_stream_conv2d_4_source_35_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_35_source_pat_fsm_17 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_35_source_ram_renable <= 0;
        _stream_conv2d_4_source_35_idle <= 1;
      end 
      if((_stream_conv2d_4_source_35_source_pat_fsm_17 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_35_source_ram_renable <= 0;
        _stream_conv2d_4_source_35_idle <= 1;
      end 
      if(_set_flag_507) begin
        _stream_conv2d_4_source_36_source_mode <= 5'b10;
        _stream_conv2d_4_source_36_source_offset <= conv2d_4_filter_page_comp_offset_buf;
      end 
      if(_set_flag_507) begin
        _source_stream_conv2d_4_source_36_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_36_pat_stride_0 <= 1;
      end 
      if(_set_flag_507) begin
        _source_stream_conv2d_4_source_36_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_36_pat_stride_1 <= cparam_conv2d_4_stream_aligned_reduce_size;
      end 
      if(_set_flag_507) begin
        _source_stream_conv2d_4_source_36_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_36_pat_stride_2 <= 0;
      end 
      if(_set_flag_507) begin
        _source_stream_conv2d_4_source_36_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_36_pat_stride_3 <= 0;
      end 
      if(_set_flag_507) begin
        _stream_conv2d_4_source_36_source_sel <= 19;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_36_source_offset_buf <= _stream_conv2d_4_source_36_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_count_0 <= _source_stream_conv2d_4_source_36_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_count_1 <= _source_stream_conv2d_4_source_36_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_count_2 <= _source_stream_conv2d_4_source_36_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_count_3 <= _source_stream_conv2d_4_source_36_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_size_buf_0 <= _source_stream_conv2d_4_source_36_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_size_buf_1 <= _source_stream_conv2d_4_source_36_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_size_buf_2 <= _source_stream_conv2d_4_source_36_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_size_buf_3 <= _source_stream_conv2d_4_source_36_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_stride_buf_0 <= _source_stream_conv2d_4_source_36_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_stride_buf_1 <= _source_stream_conv2d_4_source_36_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_stride_buf_2 <= _source_stream_conv2d_4_source_36_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_stride_buf_3 <= _source_stream_conv2d_4_source_36_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_1843 <= _stream_conv2d_4_source_36_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_36_source_pat_fsm_18 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_36_idle <= 0;
        _stream_conv2d_4_source_36_source_ram_raddr <= _stream_conv2d_4_source_36_source_pat_all_offset;
        _stream_conv2d_4_source_36_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_36_source_pat_fsm_18 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_cur_offset_0 <= _source_stream_conv2d_4_source_36_pat_cur_offset_0 + _source_stream_conv2d_4_source_36_pat_stride_buf_0;
        _source_stream_conv2d_4_source_36_pat_count_0 <= _source_stream_conv2d_4_source_36_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_36_source_pat_fsm_18 == 1) && (_source_stream_conv2d_4_source_36_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_36_pat_count_0 <= _source_stream_conv2d_4_source_36_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_36_source_pat_fsm_18 == 1) && (_source_stream_conv2d_4_source_36_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_cur_offset_1 <= _source_stream_conv2d_4_source_36_pat_cur_offset_1 + _source_stream_conv2d_4_source_36_pat_stride_buf_1;
        _source_stream_conv2d_4_source_36_pat_count_1 <= _source_stream_conv2d_4_source_36_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_36_source_pat_fsm_18 == 1) && (_source_stream_conv2d_4_source_36_pat_count_0 == 0) && (_source_stream_conv2d_4_source_36_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_36_pat_count_1 <= _source_stream_conv2d_4_source_36_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_36_source_pat_fsm_18 == 1) && ((_source_stream_conv2d_4_source_36_pat_count_0 == 0) && (_source_stream_conv2d_4_source_36_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_cur_offset_2 <= _source_stream_conv2d_4_source_36_pat_cur_offset_2 + _source_stream_conv2d_4_source_36_pat_stride_buf_2;
        _source_stream_conv2d_4_source_36_pat_count_2 <= _source_stream_conv2d_4_source_36_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_36_source_pat_fsm_18 == 1) && ((_source_stream_conv2d_4_source_36_pat_count_0 == 0) && (_source_stream_conv2d_4_source_36_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_36_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_36_pat_count_2 <= _source_stream_conv2d_4_source_36_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_36_source_pat_fsm_18 == 1) && ((_source_stream_conv2d_4_source_36_pat_count_0 == 0) && (_source_stream_conv2d_4_source_36_pat_count_1 == 0) && (_source_stream_conv2d_4_source_36_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_cur_offset_3 <= _source_stream_conv2d_4_source_36_pat_cur_offset_3 + _source_stream_conv2d_4_source_36_pat_stride_buf_3;
        _source_stream_conv2d_4_source_36_pat_count_3 <= _source_stream_conv2d_4_source_36_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_36_source_pat_fsm_18 == 1) && ((_source_stream_conv2d_4_source_36_pat_count_0 == 0) && (_source_stream_conv2d_4_source_36_pat_count_1 == 0) && (_source_stream_conv2d_4_source_36_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_36_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_36_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_36_pat_count_3 <= _source_stream_conv2d_4_source_36_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_36_source_pat_fsm_18 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_36_source_ram_renable <= 0;
        _stream_conv2d_4_source_36_idle <= 1;
      end 
      if((_stream_conv2d_4_source_36_source_pat_fsm_18 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_36_source_ram_renable <= 0;
        _stream_conv2d_4_source_36_idle <= 1;
      end 
      if(_set_flag_516) begin
        _stream_conv2d_4_source_37_source_mode <= 5'b10;
        _stream_conv2d_4_source_37_source_offset <= conv2d_4_filter_page_comp_offset_buf;
      end 
      if(_set_flag_516) begin
        _source_stream_conv2d_4_source_37_pat_size_0 <= cparam_conv2d_4_stream_reduce_size;
        _source_stream_conv2d_4_source_37_pat_stride_0 <= 1;
      end 
      if(_set_flag_516) begin
        _source_stream_conv2d_4_source_37_pat_size_1 <= conv2d_4_next_stream_num_ops;
        _source_stream_conv2d_4_source_37_pat_stride_1 <= cparam_conv2d_4_stream_aligned_reduce_size;
      end 
      if(_set_flag_516) begin
        _source_stream_conv2d_4_source_37_pat_size_2 <= 1;
        _source_stream_conv2d_4_source_37_pat_stride_2 <= 0;
      end 
      if(_set_flag_516) begin
        _source_stream_conv2d_4_source_37_pat_size_3 <= 1;
        _source_stream_conv2d_4_source_37_pat_stride_3 <= 0;
      end 
      if(_set_flag_516) begin
        _stream_conv2d_4_source_37_source_sel <= 20;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_37_source_offset_buf <= _stream_conv2d_4_source_37_source_offset;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_cur_offset_0 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_cur_offset_1 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_cur_offset_2 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_cur_offset_3 <= 0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_count_0 <= _source_stream_conv2d_4_source_37_pat_size_0 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_count_1 <= _source_stream_conv2d_4_source_37_pat_size_1 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_count_2 <= _source_stream_conv2d_4_source_37_pat_size_2 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_count_3 <= _source_stream_conv2d_4_source_37_pat_size_3 - 1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_size_buf_0 <= _source_stream_conv2d_4_source_37_pat_size_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_size_buf_1 <= _source_stream_conv2d_4_source_37_pat_size_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_size_buf_2 <= _source_stream_conv2d_4_source_37_pat_size_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_size_buf_3 <= _source_stream_conv2d_4_source_37_pat_size_3;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_stride_buf_0 <= _source_stream_conv2d_4_source_37_pat_stride_0;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_stride_buf_1 <= _source_stream_conv2d_4_source_37_pat_stride_1;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_stride_buf_2 <= _source_stream_conv2d_4_source_37_pat_stride_2;
      end 
      if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_stride_buf_3 <= _source_stream_conv2d_4_source_37_pat_stride_3;
      end 
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_busy && _stream_conv2d_4_is_root) begin
        __variable_wdata_1844 <= _stream_conv2d_4_source_37_source_ram_rdata;
      end 
      if((_stream_conv2d_4_source_37_source_pat_fsm_19 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_37_idle <= 0;
        _stream_conv2d_4_source_37_source_ram_raddr <= _stream_conv2d_4_source_37_source_pat_all_offset;
        _stream_conv2d_4_source_37_source_ram_renable <= 1;
      end 
      if((_stream_conv2d_4_source_37_source_pat_fsm_19 == 1) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_cur_offset_0 <= _source_stream_conv2d_4_source_37_pat_cur_offset_0 + _source_stream_conv2d_4_source_37_pat_stride_buf_0;
        _source_stream_conv2d_4_source_37_pat_count_0 <= _source_stream_conv2d_4_source_37_pat_count_0 - 1;
      end 
      if((_stream_conv2d_4_source_37_source_pat_fsm_19 == 1) && (_source_stream_conv2d_4_source_37_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_cur_offset_0 <= 0;
        _source_stream_conv2d_4_source_37_pat_count_0 <= _source_stream_conv2d_4_source_37_pat_size_buf_0 - 1;
      end 
      if((_stream_conv2d_4_source_37_source_pat_fsm_19 == 1) && (_source_stream_conv2d_4_source_37_pat_count_0 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_cur_offset_1 <= _source_stream_conv2d_4_source_37_pat_cur_offset_1 + _source_stream_conv2d_4_source_37_pat_stride_buf_1;
        _source_stream_conv2d_4_source_37_pat_count_1 <= _source_stream_conv2d_4_source_37_pat_count_1 - 1;
      end 
      if((_stream_conv2d_4_source_37_source_pat_fsm_19 == 1) && (_source_stream_conv2d_4_source_37_pat_count_0 == 0) && (_source_stream_conv2d_4_source_37_pat_count_1 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_cur_offset_1 <= 0;
        _source_stream_conv2d_4_source_37_pat_count_1 <= _source_stream_conv2d_4_source_37_pat_size_buf_1 - 1;
      end 
      if((_stream_conv2d_4_source_37_source_pat_fsm_19 == 1) && ((_source_stream_conv2d_4_source_37_pat_count_0 == 0) && (_source_stream_conv2d_4_source_37_pat_count_1 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_cur_offset_2 <= _source_stream_conv2d_4_source_37_pat_cur_offset_2 + _source_stream_conv2d_4_source_37_pat_stride_buf_2;
        _source_stream_conv2d_4_source_37_pat_count_2 <= _source_stream_conv2d_4_source_37_pat_count_2 - 1;
      end 
      if((_stream_conv2d_4_source_37_source_pat_fsm_19 == 1) && ((_source_stream_conv2d_4_source_37_pat_count_0 == 0) && (_source_stream_conv2d_4_source_37_pat_count_1 == 0)) && (_source_stream_conv2d_4_source_37_pat_count_2 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_cur_offset_2 <= 0;
        _source_stream_conv2d_4_source_37_pat_count_2 <= _source_stream_conv2d_4_source_37_pat_size_buf_2 - 1;
      end 
      if((_stream_conv2d_4_source_37_source_pat_fsm_19 == 1) && ((_source_stream_conv2d_4_source_37_pat_count_0 == 0) && (_source_stream_conv2d_4_source_37_pat_count_1 == 0) && (_source_stream_conv2d_4_source_37_pat_count_2 == 0)) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_cur_offset_3 <= _source_stream_conv2d_4_source_37_pat_cur_offset_3 + _source_stream_conv2d_4_source_37_pat_stride_buf_3;
        _source_stream_conv2d_4_source_37_pat_count_3 <= _source_stream_conv2d_4_source_37_pat_count_3 - 1;
      end 
      if((_stream_conv2d_4_source_37_source_pat_fsm_19 == 1) && ((_source_stream_conv2d_4_source_37_pat_count_0 == 0) && (_source_stream_conv2d_4_source_37_pat_count_1 == 0) && (_source_stream_conv2d_4_source_37_pat_count_2 == 0)) && (_source_stream_conv2d_4_source_37_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
        _source_stream_conv2d_4_source_37_pat_cur_offset_3 <= 0;
        _source_stream_conv2d_4_source_37_pat_count_3 <= _source_stream_conv2d_4_source_37_pat_size_buf_3 - 1;
      end 
      if((_stream_conv2d_4_source_37_source_pat_fsm_19 == 1) && _stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_37_source_ram_renable <= 0;
        _stream_conv2d_4_source_37_idle <= 1;
      end 
      if((_stream_conv2d_4_source_37_source_pat_fsm_19 == 2) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_source_37_source_ram_renable <= 0;
        _stream_conv2d_4_source_37_idle <= 1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_526 <= _set_flag_525;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_527 <= _tmp_526;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_528 <= _tmp_527;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_529 <= _tmp_528;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_530 <= _tmp_529;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_531 <= _tmp_530;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_532 <= _tmp_531;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_533 <= _tmp_532;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_534 <= _tmp_533;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_535 <= _tmp_534;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_536 <= _tmp_535;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_537 <= _tmp_536;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_538 <= _tmp_537;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_539 <= _tmp_538;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_540 <= _tmp_539;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_541 <= _tmp_540;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_542 <= _tmp_541;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_543 <= _tmp_542;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_544 <= _tmp_543;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_545 <= _tmp_544;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_546 <= _tmp_545;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_547 <= _tmp_546;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_548 <= _tmp_547;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_549 <= _tmp_548;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_550 <= _tmp_549;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_551 <= _tmp_550;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_552 <= _tmp_551;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_553 <= _tmp_552;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_554 <= _tmp_553;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_555 <= _tmp_554;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_556 <= _tmp_555;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_557 <= _tmp_556;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_558 <= _tmp_557;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_561 <= _tmp_560;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_562 <= _tmp_561;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_563 <= _tmp_562;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_564 <= _tmp_563;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_565 <= _tmp_564;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_566 <= _tmp_565;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_567 <= _tmp_566;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_568 <= _tmp_567;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_569 <= _tmp_568;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_570 <= _tmp_569;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_571 <= _tmp_570;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_572 <= _tmp_571;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_573 <= _tmp_572;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_574 <= _tmp_573;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_575 <= _tmp_574;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_576 <= _tmp_575;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_577 <= _tmp_576;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_578 <= _tmp_577;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_579 <= _tmp_578;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_580 <= _tmp_579;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_581 <= _tmp_580;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_582 <= _tmp_581;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_583 <= _tmp_582;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_584 <= _tmp_583;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_585 <= _tmp_584;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_586 <= _tmp_585;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_587 <= _tmp_586;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_588 <= _tmp_587;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_589 <= _tmp_588;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_590 <= _tmp_589;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_591 <= _tmp_590;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_592 <= _tmp_591;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_593 <= _tmp_592;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_594 <= conv2d_4_next_stream_num_ops;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_595 <= _tmp_594;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_596 <= _tmp_595;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_597 <= _tmp_596;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_598 <= _tmp_597;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_599 <= _tmp_598;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_600 <= _tmp_599;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_601 <= _tmp_600;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_602 <= _tmp_601;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_603 <= _tmp_602;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_604 <= _tmp_603;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_605 <= _tmp_604;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_606 <= _tmp_605;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_607 <= _tmp_606;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_608 <= _tmp_607;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_609 <= _tmp_608;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_610 <= _tmp_609;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_611 <= _tmp_610;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_612 <= _tmp_611;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_613 <= _tmp_612;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_614 <= _tmp_613;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_615 <= _tmp_614;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_616 <= _tmp_615;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_617 <= _tmp_616;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_618 <= _tmp_617;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_619 <= _tmp_618;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_620 <= _tmp_619;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_621 <= _tmp_620;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_622 <= _tmp_621;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_623 <= _tmp_622;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_624 <= _tmp_623;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_625 <= _tmp_624;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_626 <= _tmp_625;
      end 
      if(_tmp_558) begin
        _stream_conv2d_4_sink_50_sink_mode <= 5'b1;
        _stream_conv2d_4_sink_50_sink_offset <= _tmp_593;
        _stream_conv2d_4_sink_50_sink_size <= _tmp_626;
        _stream_conv2d_4_sink_50_sink_stride <= 1;
      end 
      if(_tmp_558) begin
        _stream_conv2d_4_sink_50_sink_sel <= 21;
      end 
      if(_stream_conv2d_4_sink_start && _stream_conv2d_4_sink_50_sink_mode & 5'b1 && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_sink_50_sink_offset_buf <= _stream_conv2d_4_sink_50_sink_offset;
        _stream_conv2d_4_sink_50_sink_size_buf <= _stream_conv2d_4_sink_50_sink_size;
        _stream_conv2d_4_sink_50_sink_stride_buf <= _stream_conv2d_4_sink_50_sink_stride;
      end 
      if((_stream_conv2d_4_sink_50_sink_fsm_20 == 1) && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_sink_50_sink_waddr <= _stream_conv2d_4_sink_50_sink_offset_buf - _stream_conv2d_4_sink_50_sink_stride_buf;
        _stream_conv2d_4_sink_50_sink_count <= _stream_conv2d_4_sink_50_sink_size_buf;
      end 
      if((_stream_conv2d_4_sink_50_sink_fsm_20 == 2) && stream_conv2d_4_sink_51_data && _stream_conv2d_4_stream_oready) begin
        _stream_conv2d_4_sink_50_sink_waddr <= _stream_conv2d_4_sink_50_sink_waddr + _stream_conv2d_4_sink_50_sink_stride_buf;
        _stream_conv2d_4_sink_50_sink_wdata <= stream_conv2d_4_sink_50_data;
        _stream_conv2d_4_sink_50_sink_wenable <= 1;
        _stream_conv2d_4_sink_50_sink_count <= _stream_conv2d_4_sink_50_sink_count - 1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1017 <= _stream_conv2d_4_source_start;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1018 <= _tmp_1017;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1019 <= _tmp_1018;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1020 <= _stream_conv2d_4_source_start;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1021 <= _tmp_1020;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1022 <= _tmp_1021;
      end 
      if(_stream_conv2d_4_stream_oready && _tmp_1022) begin
        __variable_wdata_1553 <= 1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1023 <= _stream_conv2d_4_source_start;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1024 <= _tmp_1023;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1025 <= _tmp_1024;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1026 <= _tmp_1025;
      end 
      if(_stream_conv2d_4_stream_oready && _tmp_1026) begin
        __variable_wdata_1553 <= 0;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1029 <= _tmp_1028;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1032 <= _tmp_1031;
      end 
      if(_stream_conv2d_4_stream_oready && _tmp_1032) begin
        __variable_wdata_1553 <= 1;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1033 <= _stream_conv2d_4_source_start;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1034 <= _tmp_1033;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1035 <= _tmp_1034;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1036 <= _tmp_1035;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1037 <= _tmp_1036;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1038 <= _tmp_1037;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1039 <= _tmp_1038;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1040 <= _tmp_1039;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1041 <= _tmp_1040;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1042 <= _tmp_1041;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1043 <= _tmp_1042;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1044 <= _tmp_1043;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1045 <= _tmp_1044;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1046 <= _tmp_1045;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1047 <= _tmp_1046;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1048 <= _tmp_1047;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1049 <= _tmp_1048;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1050 <= _tmp_1049;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1051 <= _tmp_1050;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1052 <= _tmp_1051;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1053 <= _tmp_1052;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1054 <= _tmp_1053;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1055 <= _tmp_1054;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1056 <= _tmp_1055;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1057 <= _tmp_1056;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1058 <= _tmp_1057;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1059 <= _tmp_1058;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1060 <= _tmp_1059;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1061 <= _tmp_1060;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1062 <= _tmp_1061;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1063 <= _tmp_1062;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1064 <= _tmp_1063;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1065 <= _tmp_1064;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1066 <= _stream_conv2d_4_source_stop;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1067 <= _tmp_1066;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1068 <= _tmp_1067;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1069 <= _tmp_1068;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1070 <= _tmp_1069;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1071 <= _tmp_1070;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1072 <= _tmp_1071;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1073 <= _tmp_1072;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1074 <= _tmp_1073;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1075 <= _tmp_1074;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1076 <= _tmp_1075;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1077 <= _tmp_1076;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1078 <= _tmp_1077;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1079 <= _tmp_1078;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1080 <= _tmp_1079;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1081 <= _tmp_1080;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1082 <= _tmp_1081;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1083 <= _tmp_1082;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1084 <= _tmp_1083;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1085 <= _tmp_1084;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1086 <= _tmp_1085;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1087 <= _tmp_1086;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1088 <= _tmp_1087;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1089 <= _tmp_1088;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1090 <= _tmp_1089;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1091 <= _tmp_1090;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1092 <= _tmp_1091;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1093 <= _tmp_1092;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1094 <= _tmp_1093;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1095 <= _tmp_1094;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1096 <= _tmp_1095;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1097 <= _tmp_1096;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1098 <= _tmp_1097;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1099 <= _stream_conv2d_4_source_busy;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1100 <= _tmp_1099;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1101 <= _tmp_1100;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1102 <= _tmp_1101;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1103 <= _tmp_1102;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1104 <= _tmp_1103;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1105 <= _tmp_1104;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1106 <= _tmp_1105;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1107 <= _tmp_1106;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1108 <= _tmp_1107;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1109 <= _tmp_1108;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1110 <= _tmp_1109;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1111 <= _tmp_1110;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1112 <= _tmp_1111;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1113 <= _tmp_1112;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1114 <= _tmp_1113;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1115 <= _tmp_1114;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1116 <= _tmp_1115;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1117 <= _tmp_1116;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1118 <= _tmp_1117;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1119 <= _tmp_1118;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1120 <= _tmp_1119;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1121 <= _tmp_1120;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1122 <= _tmp_1121;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1123 <= _tmp_1122;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1124 <= _tmp_1123;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1125 <= _tmp_1124;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1126 <= _tmp_1125;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1127 <= _tmp_1126;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1128 <= _tmp_1127;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1129 <= _tmp_1128;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1130 <= _tmp_1129;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1131 <= _tmp_1130;
      end 
      if(_stream_conv2d_4_stream_oready) begin
        _tmp_1132 <= _stream_conv2d_4_sink_busy;
      end 
      if(!_stream_conv2d_4_sink_busy && _tmp_1132) begin
        _stream_conv2d_4_busy_reg <= 0;
      end 
      if(_stream_conv2d_4_source_busy) begin
        _stream_conv2d_4_busy_reg <= 1;
      end 
    end
  end

  localparam _stream_conv2d_4_fsm_1 = 1;
  localparam _stream_conv2d_4_fsm_2 = 2;
  localparam _stream_conv2d_4_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_fsm <= _stream_conv2d_4_fsm_init;
      _stream_conv2d_4_source_start <= 0;
      _stream_conv2d_4_source_busy <= 0;
      _stream_conv2d_4_stream_ivalid <= 0;
    end else begin
      if(_stream_conv2d_4_stream_oready && _tmp_1019) begin
        _stream_conv2d_4_stream_ivalid <= 1;
      end 
      if(_stream_conv2d_4_stream_oready && _tmp_1029) begin
        _stream_conv2d_4_stream_ivalid <= 0;
      end 
      case(_stream_conv2d_4_fsm)
        _stream_conv2d_4_fsm_init: begin
          if(_stream_conv2d_4_run_flag) begin
            _stream_conv2d_4_source_start <= 1;
          end 
          if(_stream_conv2d_4_run_flag) begin
            _stream_conv2d_4_fsm <= _stream_conv2d_4_fsm_1;
          end 
        end
        _stream_conv2d_4_fsm_1: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_start <= 0;
            _stream_conv2d_4_source_busy <= 1;
          end 
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_fsm <= _stream_conv2d_4_fsm_2;
          end 
        end
        _stream_conv2d_4_fsm_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_fsm <= _stream_conv2d_4_fsm_3;
          end 
        end
        _stream_conv2d_4_fsm_3: begin
          if(_stream_conv2d_4_stream_oready && (_stream_conv2d_4_source_11_idle && _stream_conv2d_4_source_13_idle && _stream_conv2d_4_source_15_idle && _stream_conv2d_4_source_20_idle && _stream_conv2d_4_source_21_idle && _stream_conv2d_4_source_22_idle && _stream_conv2d_4_source_23_idle && _stream_conv2d_4_source_24_idle && _stream_conv2d_4_source_25_idle && _stream_conv2d_4_source_26_idle && _stream_conv2d_4_source_27_idle && _stream_conv2d_4_source_28_idle && _stream_conv2d_4_source_29_idle && _stream_conv2d_4_source_30_idle && _stream_conv2d_4_source_31_idle && _stream_conv2d_4_source_32_idle && _stream_conv2d_4_source_33_idle && _stream_conv2d_4_source_34_idle && _stream_conv2d_4_source_35_idle && _stream_conv2d_4_source_36_idle && _stream_conv2d_4_source_37_idle && _stream_conv2d_4_source_7_idle && _stream_conv2d_4_source_9_idle && (_stream_conv2d_4_fsm == 3))) begin
            _stream_conv2d_4_source_busy <= 0;
          end 
          if(_stream_conv2d_4_stream_oready && (_stream_conv2d_4_source_11_idle && _stream_conv2d_4_source_13_idle && _stream_conv2d_4_source_15_idle && _stream_conv2d_4_source_20_idle && _stream_conv2d_4_source_21_idle && _stream_conv2d_4_source_22_idle && _stream_conv2d_4_source_23_idle && _stream_conv2d_4_source_24_idle && _stream_conv2d_4_source_25_idle && _stream_conv2d_4_source_26_idle && _stream_conv2d_4_source_27_idle && _stream_conv2d_4_source_28_idle && _stream_conv2d_4_source_29_idle && _stream_conv2d_4_source_30_idle && _stream_conv2d_4_source_31_idle && _stream_conv2d_4_source_32_idle && _stream_conv2d_4_source_33_idle && _stream_conv2d_4_source_34_idle && _stream_conv2d_4_source_35_idle && _stream_conv2d_4_source_36_idle && _stream_conv2d_4_source_37_idle && _stream_conv2d_4_source_7_idle && _stream_conv2d_4_source_9_idle && (_stream_conv2d_4_fsm == 3)) && _stream_conv2d_4_run_flag) begin
            _stream_conv2d_4_source_start <= 1;
          end 
          if(_stream_conv2d_4_stream_oready && (_stream_conv2d_4_source_11_idle && _stream_conv2d_4_source_13_idle && _stream_conv2d_4_source_15_idle && _stream_conv2d_4_source_20_idle && _stream_conv2d_4_source_21_idle && _stream_conv2d_4_source_22_idle && _stream_conv2d_4_source_23_idle && _stream_conv2d_4_source_24_idle && _stream_conv2d_4_source_25_idle && _stream_conv2d_4_source_26_idle && _stream_conv2d_4_source_27_idle && _stream_conv2d_4_source_28_idle && _stream_conv2d_4_source_29_idle && _stream_conv2d_4_source_30_idle && _stream_conv2d_4_source_31_idle && _stream_conv2d_4_source_32_idle && _stream_conv2d_4_source_33_idle && _stream_conv2d_4_source_34_idle && _stream_conv2d_4_source_35_idle && _stream_conv2d_4_source_36_idle && _stream_conv2d_4_source_37_idle && _stream_conv2d_4_source_7_idle && _stream_conv2d_4_source_9_idle && (_stream_conv2d_4_fsm == 3))) begin
            _stream_conv2d_4_fsm <= _stream_conv2d_4_fsm_init;
          end 
          if(_stream_conv2d_4_stream_oready && (_stream_conv2d_4_source_11_idle && _stream_conv2d_4_source_13_idle && _stream_conv2d_4_source_15_idle && _stream_conv2d_4_source_20_idle && _stream_conv2d_4_source_21_idle && _stream_conv2d_4_source_22_idle && _stream_conv2d_4_source_23_idle && _stream_conv2d_4_source_24_idle && _stream_conv2d_4_source_25_idle && _stream_conv2d_4_source_26_idle && _stream_conv2d_4_source_27_idle && _stream_conv2d_4_source_28_idle && _stream_conv2d_4_source_29_idle && _stream_conv2d_4_source_30_idle && _stream_conv2d_4_source_31_idle && _stream_conv2d_4_source_32_idle && _stream_conv2d_4_source_33_idle && _stream_conv2d_4_source_34_idle && _stream_conv2d_4_source_35_idle && _stream_conv2d_4_source_36_idle && _stream_conv2d_4_source_37_idle && _stream_conv2d_4_source_7_idle && _stream_conv2d_4_source_9_idle && (_stream_conv2d_4_fsm == 3)) && _stream_conv2d_4_run_flag) begin
            _stream_conv2d_4_fsm <= _stream_conv2d_4_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _stream_max_pool_serial_6_source_1_source_ram_renable <= 0;
      _stream_max_pool_serial_6_source_1_source_fifo_deq <= 0;
      _stream_max_pool_serial_6_source_1_idle <= 1;
      _stream_max_pool_serial_6_sink_5_sink_wenable <= 0;
      _stream_max_pool_serial_6_sink_5_sink_fifo_enq <= 0;
      _stream_max_pool_serial_6_sink_6_sink_wenable <= 0;
      _stream_max_pool_serial_6_sink_6_sink_fifo_enq <= 0;
      __stream_max_pool_serial_6_stream_ivalid_1 <= 0;
      __stream_max_pool_serial_6_stream_ivalid_2 <= 0;
      __stream_max_pool_serial_6_stream_ivalid_3 <= 0;
      __stream_max_pool_serial_6_stream_ivalid_4 <= 0;
      __stream_max_pool_serial_6_stream_ivalid_5 <= 0;
      _counter_data_2141 <= 1'sd0;
      _counter_count_2141 <= 1'sd0;
      __delay_data_2394__variable_2139 <= 0;
      __delay_data_2395_reinterpretcast_2149 <= 0;
      __delay_data_2397__variable_2140 <= 0;
      __delay_data_2400__variable_2137 <= 0;
      _pointer_data_2144 <= 0;
      __delay_data_2396__delay_2395_reinterpretcast_2149 <= 0;
      __delay_data_2398__delay_2397__variable_2140 <= 0;
      __delay_data_2401__delay_2400__variable_2137 <= 0;
      _cond_data_2151 <= 0;
      __delay_data_2399__delay_2398__delay_2397__variable_2140 <= 0;
      __delay_data_2402__delay_2401__delay_2400__variable_2137 <= 0;
      _stream_max_pool_serial_6_parameter_0_next_parameter_data <= 0;
      __variable_wdata_2137 <= 0;
      _stream_max_pool_serial_6_parameter_2_next_parameter_data <= 0;
      __variable_wdata_2139 <= 0;
      _stream_max_pool_serial_6_source_1_source_mode <= 5'b0;
      _stream_max_pool_serial_6_source_1_source_offset <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_size_0 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_stride_0 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_size_1 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_stride_1 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_size_2 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_stride_2 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_size_3 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_stride_3 <= 0;
      _stream_max_pool_serial_6_source_1_source_sel <= 0;
      _stream_max_pool_serial_6_source_1_source_offset_buf <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_cur_offset_0 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_cur_offset_1 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_cur_offset_2 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_cur_offset_3 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_count_0 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_count_1 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_count_2 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_count_3 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_size_buf_0 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_size_buf_1 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_size_buf_2 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_size_buf_3 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_stride_buf_0 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_stride_buf_1 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_stride_buf_2 <= 0;
      _source_stream_max_pool_serial_6_source_1_pat_stride_buf_3 <= 0;
      __variable_wdata_2138 <= 0;
      _stream_max_pool_serial_6_source_1_source_ram_raddr <= 0;
      _tmp_1210 <= 0;
      _tmp_1211 <= 0;
      _tmp_1212 <= 0;
      _tmp_1213 <= 0;
      _tmp_1214 <= 0;
      _tmp_1215 <= 0;
      _tmp_1216 <= 0;
      _tmp_1219 <= 0;
      _tmp_1220 <= 0;
      _tmp_1221 <= 0;
      _tmp_1222 <= 0;
      _tmp_1223 <= 0;
      _tmp_1224 <= 0;
      _tmp_1225 <= 0;
      _tmp_1226 <= 0;
      _tmp_1227 <= 0;
      _tmp_1228 <= 0;
      _tmp_1229 <= 0;
      _tmp_1230 <= 0;
      _tmp_1231 <= 0;
      _tmp_1232 <= 0;
      _stream_max_pool_serial_6_sink_5_sink_mode <= 5'b0;
      _stream_max_pool_serial_6_sink_5_sink_offset <= 0;
      _stream_max_pool_serial_6_sink_5_sink_size <= 0;
      _stream_max_pool_serial_6_sink_5_sink_stride <= 0;
      _stream_max_pool_serial_6_sink_5_sink_sel <= 0;
      _stream_max_pool_serial_6_sink_5_sink_offset_buf <= 0;
      _stream_max_pool_serial_6_sink_5_sink_size_buf <= 0;
      _stream_max_pool_serial_6_sink_5_sink_stride_buf <= 0;
      _stream_max_pool_serial_6_sink_5_sink_waddr <= 0;
      _stream_max_pool_serial_6_sink_5_sink_count <= 0;
      _stream_max_pool_serial_6_sink_5_sink_wdata <= 0;
      _tmp_1255 <= 0;
      _tmp_1256 <= 0;
      _tmp_1257 <= 0;
      _tmp_1258 <= 0;
      _tmp_1259 <= 0;
      _tmp_1260 <= 0;
      __variable_wdata_2140 <= 0;
      _tmp_1261 <= 0;
      _tmp_1262 <= 0;
      _tmp_1263 <= 0;
      _tmp_1264 <= 0;
      _tmp_1267 <= 0;
      _tmp_1270 <= 0;
      _tmp_1271 <= 0;
      _tmp_1272 <= 0;
      _tmp_1273 <= 0;
      _tmp_1274 <= 0;
      _tmp_1275 <= 0;
      _tmp_1276 <= 0;
      _tmp_1277 <= 0;
      _tmp_1278 <= 0;
      _tmp_1279 <= 0;
      _tmp_1280 <= 0;
      _tmp_1281 <= 0;
      _tmp_1282 <= 0;
      _tmp_1283 <= 0;
      _tmp_1284 <= 0;
      _tmp_1285 <= 0;
      _tmp_1286 <= 0;
      _tmp_1287 <= 0;
      _tmp_1288 <= 0;
      _tmp_1289 <= 0;
      _tmp_1290 <= 0;
      _tmp_1291 <= 0;
      _tmp_1292 <= 0;
      _stream_max_pool_serial_6_busy_reg <= 0;
    end else begin
      if(_stream_max_pool_serial_6_stream_oready) begin
        _stream_max_pool_serial_6_source_1_source_ram_renable <= 0;
        _stream_max_pool_serial_6_source_1_source_fifo_deq <= 0;
      end 
      _stream_max_pool_serial_6_source_1_idle <= _stream_max_pool_serial_6_source_1_idle;
      if(_stream_max_pool_serial_6_stream_oready) begin
        _stream_max_pool_serial_6_sink_5_sink_wenable <= 0;
        _stream_max_pool_serial_6_sink_5_sink_fifo_enq <= 0;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _stream_max_pool_serial_6_sink_6_sink_wenable <= 0;
        _stream_max_pool_serial_6_sink_6_sink_fifo_enq <= 0;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        __stream_max_pool_serial_6_stream_ivalid_1 <= _stream_max_pool_serial_6_stream_ivalid;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        __stream_max_pool_serial_6_stream_ivalid_2 <= __stream_max_pool_serial_6_stream_ivalid_1;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        __stream_max_pool_serial_6_stream_ivalid_3 <= __stream_max_pool_serial_6_stream_ivalid_2;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        __stream_max_pool_serial_6_stream_ivalid_4 <= __stream_max_pool_serial_6_stream_ivalid_3;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        __stream_max_pool_serial_6_stream_ivalid_5 <= __stream_max_pool_serial_6_stream_ivalid_4;
      end 
      if(_stream_max_pool_serial_6_stream_ivalid && _stream_max_pool_serial_6_stream_oready && _counter_reset_cond_2141) begin
        _counter_data_2141 <= 1'sd0;
      end 
      if(_stream_max_pool_serial_6_stream_ivalid && _stream_max_pool_serial_6_stream_oready) begin
        _counter_data_2141 <= _counter_current_count_2141;
      end 
      if(_stream_max_pool_serial_6_stream_ivalid && _stream_max_pool_serial_6_stream_oready) begin
        _counter_count_2141 <= (_counter_current_count_2141 >= stream_max_pool_serial_6_parameter_0_data - 2'sd1)? _counter_current_count_2141 + 2'sd1 - stream_max_pool_serial_6_parameter_0_data : _counter_current_count_2141 + 2'sd1;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        __delay_data_2394__variable_2139 <= stream_max_pool_serial_6_parameter_2_data;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        __delay_data_2395_reinterpretcast_2149 <= _reinterpretcast_data_2149;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        __delay_data_2397__variable_2140 <= stream_max_pool_serial_6__reduce_reset_data;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        __delay_data_2400__variable_2137 <= stream_max_pool_serial_6_parameter_0_data;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _pointer_data_2144 <= __delay_data_2394__variable_2139[_counter_data_2141];
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        __delay_data_2396__delay_2395_reinterpretcast_2149 <= __delay_data_2395_reinterpretcast_2149;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        __delay_data_2398__delay_2397__variable_2140 <= __delay_data_2397__variable_2140;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        __delay_data_2401__delay_2400__variable_2137 <= __delay_data_2400__variable_2137;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _cond_data_2151 <= (_pointer_data_2144)? -17'sd32768 : __delay_data_2396__delay_2395_reinterpretcast_2149;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        __delay_data_2399__delay_2398__delay_2397__variable_2140 <= __delay_data_2398__delay_2397__variable_2140;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        __delay_data_2402__delay_2401__delay_2400__variable_2137 <= __delay_data_2401__delay_2400__variable_2137;
      end 
      if(_set_flag_1198) begin
        _stream_max_pool_serial_6_parameter_0_next_parameter_data <= 4;
      end 
      if(_stream_max_pool_serial_6_source_start) begin
        __variable_wdata_2137 <= _stream_max_pool_serial_6_parameter_0_next_parameter_data;
      end 
      if(_set_flag_1199) begin
        _stream_max_pool_serial_6_parameter_2_next_parameter_data <= max_pool_serial_6_stream_pad_masks;
      end 
      if(_stream_max_pool_serial_6_source_start) begin
        __variable_wdata_2139 <= _stream_max_pool_serial_6_parameter_2_next_parameter_data;
      end 
      if(_set_flag_1200) begin
        _stream_max_pool_serial_6_source_1_source_mode <= 5'b10;
        _stream_max_pool_serial_6_source_1_source_offset <= max_pool_serial_6_stream_act_local + max_pool_serial_6_act_page_comp_offset_buf;
      end 
      if(_set_flag_1200) begin
        _source_stream_max_pool_serial_6_source_1_pat_size_0 <= 2;
        _source_stream_max_pool_serial_6_source_1_pat_stride_0 <= cparam_max_pool_serial_6_act_read_block;
      end 
      if(_set_flag_1200) begin
        _source_stream_max_pool_serial_6_source_1_pat_size_1 <= 2;
        _source_stream_max_pool_serial_6_source_1_pat_stride_1 <= cparam_max_pool_serial_6_act_read_size;
      end 
      if(_set_flag_1200) begin
        _source_stream_max_pool_serial_6_source_1_pat_size_2 <= cparam_max_pool_serial_6_stream_size;
        _source_stream_max_pool_serial_6_source_1_pat_stride_2 <= 1;
      end 
      if(_set_flag_1200) begin
        _source_stream_max_pool_serial_6_source_1_pat_size_3 <= 1;
        _source_stream_max_pool_serial_6_source_1_pat_stride_3 <= 0;
      end 
      if(_set_flag_1200) begin
        _stream_max_pool_serial_6_source_1_source_sel <= 1;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _stream_max_pool_serial_6_source_1_source_offset_buf <= _stream_max_pool_serial_6_source_1_source_offset;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_cur_offset_0 <= 0;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_cur_offset_1 <= 0;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_cur_offset_2 <= 0;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_cur_offset_3 <= 0;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_count_0 <= _source_stream_max_pool_serial_6_source_1_pat_size_0 - 1;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_count_1 <= _source_stream_max_pool_serial_6_source_1_pat_size_1 - 1;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_count_2 <= _source_stream_max_pool_serial_6_source_1_pat_size_2 - 1;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_count_3 <= _source_stream_max_pool_serial_6_source_1_pat_size_3 - 1;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_size_buf_0 <= _source_stream_max_pool_serial_6_source_1_pat_size_0;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_size_buf_1 <= _source_stream_max_pool_serial_6_source_1_pat_size_1;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_size_buf_2 <= _source_stream_max_pool_serial_6_source_1_pat_size_2;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_size_buf_3 <= _source_stream_max_pool_serial_6_source_1_pat_size_3;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_stride_buf_0 <= _source_stream_max_pool_serial_6_source_1_pat_stride_0;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_stride_buf_1 <= _source_stream_max_pool_serial_6_source_1_pat_stride_1;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_stride_buf_2 <= _source_stream_max_pool_serial_6_source_1_pat_stride_2;
      end 
      if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_stride_buf_3 <= _source_stream_max_pool_serial_6_source_1_pat_stride_3;
      end 
      if(_stream_max_pool_serial_6_stream_oready && _stream_max_pool_serial_6_source_busy && _stream_max_pool_serial_6_is_root) begin
        __variable_wdata_2138 <= _stream_max_pool_serial_6_source_1_source_ram_rdata;
      end 
      if((_stream_max_pool_serial_6_source_1_source_pat_fsm_0 == 1) && _stream_max_pool_serial_6_stream_oready) begin
        _stream_max_pool_serial_6_source_1_idle <= 0;
        _stream_max_pool_serial_6_source_1_source_ram_raddr <= _stream_max_pool_serial_6_source_1_source_pat_all_offset;
        _stream_max_pool_serial_6_source_1_source_ram_renable <= 1;
      end 
      if((_stream_max_pool_serial_6_source_1_source_pat_fsm_0 == 1) && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_cur_offset_0 <= _source_stream_max_pool_serial_6_source_1_pat_cur_offset_0 + _source_stream_max_pool_serial_6_source_1_pat_stride_buf_0;
        _source_stream_max_pool_serial_6_source_1_pat_count_0 <= _source_stream_max_pool_serial_6_source_1_pat_count_0 - 1;
      end 
      if((_stream_max_pool_serial_6_source_1_source_pat_fsm_0 == 1) && (_source_stream_max_pool_serial_6_source_1_pat_count_0 == 0) && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_cur_offset_0 <= 0;
        _source_stream_max_pool_serial_6_source_1_pat_count_0 <= _source_stream_max_pool_serial_6_source_1_pat_size_buf_0 - 1;
      end 
      if((_stream_max_pool_serial_6_source_1_source_pat_fsm_0 == 1) && (_source_stream_max_pool_serial_6_source_1_pat_count_0 == 0) && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_cur_offset_1 <= _source_stream_max_pool_serial_6_source_1_pat_cur_offset_1 + _source_stream_max_pool_serial_6_source_1_pat_stride_buf_1;
        _source_stream_max_pool_serial_6_source_1_pat_count_1 <= _source_stream_max_pool_serial_6_source_1_pat_count_1 - 1;
      end 
      if((_stream_max_pool_serial_6_source_1_source_pat_fsm_0 == 1) && (_source_stream_max_pool_serial_6_source_1_pat_count_0 == 0) && (_source_stream_max_pool_serial_6_source_1_pat_count_1 == 0) && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_cur_offset_1 <= 0;
        _source_stream_max_pool_serial_6_source_1_pat_count_1 <= _source_stream_max_pool_serial_6_source_1_pat_size_buf_1 - 1;
      end 
      if((_stream_max_pool_serial_6_source_1_source_pat_fsm_0 == 1) && ((_source_stream_max_pool_serial_6_source_1_pat_count_0 == 0) && (_source_stream_max_pool_serial_6_source_1_pat_count_1 == 0)) && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_cur_offset_2 <= _source_stream_max_pool_serial_6_source_1_pat_cur_offset_2 + _source_stream_max_pool_serial_6_source_1_pat_stride_buf_2;
        _source_stream_max_pool_serial_6_source_1_pat_count_2 <= _source_stream_max_pool_serial_6_source_1_pat_count_2 - 1;
      end 
      if((_stream_max_pool_serial_6_source_1_source_pat_fsm_0 == 1) && ((_source_stream_max_pool_serial_6_source_1_pat_count_0 == 0) && (_source_stream_max_pool_serial_6_source_1_pat_count_1 == 0)) && (_source_stream_max_pool_serial_6_source_1_pat_count_2 == 0) && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_cur_offset_2 <= 0;
        _source_stream_max_pool_serial_6_source_1_pat_count_2 <= _source_stream_max_pool_serial_6_source_1_pat_size_buf_2 - 1;
      end 
      if((_stream_max_pool_serial_6_source_1_source_pat_fsm_0 == 1) && ((_source_stream_max_pool_serial_6_source_1_pat_count_0 == 0) && (_source_stream_max_pool_serial_6_source_1_pat_count_1 == 0) && (_source_stream_max_pool_serial_6_source_1_pat_count_2 == 0)) && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_cur_offset_3 <= _source_stream_max_pool_serial_6_source_1_pat_cur_offset_3 + _source_stream_max_pool_serial_6_source_1_pat_stride_buf_3;
        _source_stream_max_pool_serial_6_source_1_pat_count_3 <= _source_stream_max_pool_serial_6_source_1_pat_count_3 - 1;
      end 
      if((_stream_max_pool_serial_6_source_1_source_pat_fsm_0 == 1) && ((_source_stream_max_pool_serial_6_source_1_pat_count_0 == 0) && (_source_stream_max_pool_serial_6_source_1_pat_count_1 == 0) && (_source_stream_max_pool_serial_6_source_1_pat_count_2 == 0)) && (_source_stream_max_pool_serial_6_source_1_pat_count_3 == 0) && _stream_max_pool_serial_6_stream_oready) begin
        _source_stream_max_pool_serial_6_source_1_pat_cur_offset_3 <= 0;
        _source_stream_max_pool_serial_6_source_1_pat_count_3 <= _source_stream_max_pool_serial_6_source_1_pat_size_buf_3 - 1;
      end 
      if((_stream_max_pool_serial_6_source_1_source_pat_fsm_0 == 1) && _stream_max_pool_serial_6_source_stop && _stream_max_pool_serial_6_stream_oready) begin
        _stream_max_pool_serial_6_source_1_source_ram_renable <= 0;
        _stream_max_pool_serial_6_source_1_idle <= 1;
      end 
      if((_stream_max_pool_serial_6_source_1_source_pat_fsm_0 == 2) && _stream_max_pool_serial_6_stream_oready) begin
        _stream_max_pool_serial_6_source_1_source_ram_renable <= 0;
        _stream_max_pool_serial_6_source_1_idle <= 1;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1210 <= _set_flag_1209;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1211 <= _tmp_1210;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1212 <= _tmp_1211;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1213 <= _tmp_1212;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1214 <= _tmp_1213;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1215 <= _tmp_1214;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1216 <= _tmp_1215;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1219 <= _tmp_1218;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1220 <= _tmp_1219;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1221 <= _tmp_1220;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1222 <= _tmp_1221;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1223 <= _tmp_1222;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1224 <= _tmp_1223;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1225 <= _tmp_1224;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1226 <= cparam_max_pool_serial_6_stream_size;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1227 <= _tmp_1226;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1228 <= _tmp_1227;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1229 <= _tmp_1228;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1230 <= _tmp_1229;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1231 <= _tmp_1230;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1232 <= _tmp_1231;
      end 
      if(_tmp_1216) begin
        _stream_max_pool_serial_6_sink_5_sink_mode <= 5'b1;
        _stream_max_pool_serial_6_sink_5_sink_offset <= _tmp_1225;
        _stream_max_pool_serial_6_sink_5_sink_size <= _tmp_1232;
        _stream_max_pool_serial_6_sink_5_sink_stride <= 1;
      end 
      if(_tmp_1216) begin
        _stream_max_pool_serial_6_sink_5_sink_sel <= 2;
      end 
      if(_stream_max_pool_serial_6_sink_start && _stream_max_pool_serial_6_sink_5_sink_mode & 5'b1 && _stream_max_pool_serial_6_stream_oready) begin
        _stream_max_pool_serial_6_sink_5_sink_offset_buf <= _stream_max_pool_serial_6_sink_5_sink_offset;
        _stream_max_pool_serial_6_sink_5_sink_size_buf <= _stream_max_pool_serial_6_sink_5_sink_size;
        _stream_max_pool_serial_6_sink_5_sink_stride_buf <= _stream_max_pool_serial_6_sink_5_sink_stride;
      end 
      if((_stream_max_pool_serial_6_sink_5_sink_fsm_1 == 1) && _stream_max_pool_serial_6_stream_oready) begin
        _stream_max_pool_serial_6_sink_5_sink_waddr <= _stream_max_pool_serial_6_sink_5_sink_offset_buf - _stream_max_pool_serial_6_sink_5_sink_stride_buf;
        _stream_max_pool_serial_6_sink_5_sink_count <= _stream_max_pool_serial_6_sink_5_sink_size_buf;
      end 
      if((_stream_max_pool_serial_6_sink_5_sink_fsm_1 == 2) && stream_max_pool_serial_6_sink_6_data && _stream_max_pool_serial_6_stream_oready) begin
        _stream_max_pool_serial_6_sink_5_sink_waddr <= _stream_max_pool_serial_6_sink_5_sink_waddr + _stream_max_pool_serial_6_sink_5_sink_stride_buf;
        _stream_max_pool_serial_6_sink_5_sink_wdata <= stream_max_pool_serial_6_sink_5_data;
        _stream_max_pool_serial_6_sink_5_sink_wenable <= 1;
        _stream_max_pool_serial_6_sink_5_sink_count <= _stream_max_pool_serial_6_sink_5_sink_count - 1;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1255 <= _stream_max_pool_serial_6_source_start;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1256 <= _tmp_1255;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1257 <= _tmp_1256;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1258 <= _stream_max_pool_serial_6_source_start;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1259 <= _tmp_1258;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1260 <= _tmp_1259;
      end 
      if(_stream_max_pool_serial_6_stream_oready && _tmp_1260) begin
        __variable_wdata_2140 <= 1;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1261 <= _stream_max_pool_serial_6_source_start;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1262 <= _tmp_1261;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1263 <= _tmp_1262;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1264 <= _tmp_1263;
      end 
      if(_stream_max_pool_serial_6_stream_oready && _tmp_1264) begin
        __variable_wdata_2140 <= 0;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1267 <= _tmp_1266;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1270 <= _tmp_1269;
      end 
      if(_stream_max_pool_serial_6_stream_oready && _tmp_1270) begin
        __variable_wdata_2140 <= 1;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1271 <= _stream_max_pool_serial_6_source_start;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1272 <= _tmp_1271;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1273 <= _tmp_1272;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1274 <= _tmp_1273;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1275 <= _tmp_1274;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1276 <= _tmp_1275;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1277 <= _tmp_1276;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1278 <= _stream_max_pool_serial_6_source_stop;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1279 <= _tmp_1278;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1280 <= _tmp_1279;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1281 <= _tmp_1280;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1282 <= _tmp_1281;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1283 <= _tmp_1282;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1284 <= _tmp_1283;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1285 <= _stream_max_pool_serial_6_source_busy;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1286 <= _tmp_1285;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1287 <= _tmp_1286;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1288 <= _tmp_1287;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1289 <= _tmp_1288;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1290 <= _tmp_1289;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1291 <= _tmp_1290;
      end 
      if(_stream_max_pool_serial_6_stream_oready) begin
        _tmp_1292 <= _stream_max_pool_serial_6_sink_busy;
      end 
      if(!_stream_max_pool_serial_6_sink_busy && _tmp_1292) begin
        _stream_max_pool_serial_6_busy_reg <= 0;
      end 
      if(_stream_max_pool_serial_6_source_busy) begin
        _stream_max_pool_serial_6_busy_reg <= 1;
      end 
    end
  end

  localparam _stream_max_pool_serial_6_fsm_1 = 1;
  localparam _stream_max_pool_serial_6_fsm_2 = 2;
  localparam _stream_max_pool_serial_6_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_max_pool_serial_6_fsm <= _stream_max_pool_serial_6_fsm_init;
      _stream_max_pool_serial_6_source_start <= 0;
      _stream_max_pool_serial_6_source_busy <= 0;
      _stream_max_pool_serial_6_stream_ivalid <= 0;
    end else begin
      if(_stream_max_pool_serial_6_stream_oready && _tmp_1257) begin
        _stream_max_pool_serial_6_stream_ivalid <= 1;
      end 
      if(_stream_max_pool_serial_6_stream_oready && _tmp_1267) begin
        _stream_max_pool_serial_6_stream_ivalid <= 0;
      end 
      case(_stream_max_pool_serial_6_fsm)
        _stream_max_pool_serial_6_fsm_init: begin
          if(_stream_max_pool_serial_6_run_flag) begin
            _stream_max_pool_serial_6_source_start <= 1;
          end 
          if(_stream_max_pool_serial_6_run_flag) begin
            _stream_max_pool_serial_6_fsm <= _stream_max_pool_serial_6_fsm_1;
          end 
        end
        _stream_max_pool_serial_6_fsm_1: begin
          if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_stream_oready) begin
            _stream_max_pool_serial_6_source_start <= 0;
            _stream_max_pool_serial_6_source_busy <= 1;
          end 
          if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_stream_oready) begin
            _stream_max_pool_serial_6_fsm <= _stream_max_pool_serial_6_fsm_2;
          end 
        end
        _stream_max_pool_serial_6_fsm_2: begin
          if(_stream_max_pool_serial_6_stream_oready) begin
            _stream_max_pool_serial_6_fsm <= _stream_max_pool_serial_6_fsm_3;
          end 
        end
        _stream_max_pool_serial_6_fsm_3: begin
          if(_stream_max_pool_serial_6_stream_oready && (_stream_max_pool_serial_6_source_1_idle && (_stream_max_pool_serial_6_fsm == 3))) begin
            _stream_max_pool_serial_6_source_busy <= 0;
          end 
          if(_stream_max_pool_serial_6_stream_oready && (_stream_max_pool_serial_6_source_1_idle && (_stream_max_pool_serial_6_fsm == 3)) && _stream_max_pool_serial_6_run_flag) begin
            _stream_max_pool_serial_6_source_start <= 1;
          end 
          if(_stream_max_pool_serial_6_stream_oready && (_stream_max_pool_serial_6_source_1_idle && (_stream_max_pool_serial_6_fsm == 3))) begin
            _stream_max_pool_serial_6_fsm <= _stream_max_pool_serial_6_fsm_init;
          end 
          if(_stream_max_pool_serial_6_stream_oready && (_stream_max_pool_serial_6_source_1_idle && (_stream_max_pool_serial_6_fsm == 3)) && _stream_max_pool_serial_6_run_flag) begin
            _stream_max_pool_serial_6_fsm <= _stream_max_pool_serial_6_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _stream_matmul_11_source_7_source_ram_renable <= 0;
      _stream_matmul_11_source_7_source_fifo_deq <= 0;
      _stream_matmul_11_source_7_idle <= 1;
      _stream_matmul_11_source_9_source_ram_renable <= 0;
      _stream_matmul_11_source_9_source_fifo_deq <= 0;
      _stream_matmul_11_source_9_idle <= 1;
      _stream_matmul_11_source_11_source_ram_renable <= 0;
      _stream_matmul_11_source_11_source_fifo_deq <= 0;
      _stream_matmul_11_source_11_idle <= 1;
      _stream_matmul_11_source_13_source_ram_renable <= 0;
      _stream_matmul_11_source_13_source_fifo_deq <= 0;
      _stream_matmul_11_source_13_idle <= 1;
      _stream_matmul_11_source_15_source_ram_renable <= 0;
      _stream_matmul_11_source_15_source_fifo_deq <= 0;
      _stream_matmul_11_source_15_idle <= 1;
      _stream_matmul_11_source_20_source_ram_renable <= 0;
      _stream_matmul_11_source_20_source_fifo_deq <= 0;
      _stream_matmul_11_source_20_idle <= 1;
      _stream_matmul_11_source_21_source_ram_renable <= 0;
      _stream_matmul_11_source_21_source_fifo_deq <= 0;
      _stream_matmul_11_source_21_idle <= 1;
      _stream_matmul_11_sink_26_sink_wenable <= 0;
      _stream_matmul_11_sink_26_sink_fifo_enq <= 0;
      _stream_matmul_11_sink_27_sink_wenable <= 0;
      _stream_matmul_11_sink_27_sink_fifo_enq <= 0;
      __stream_matmul_11_stream_ivalid_1 <= 0;
      __stream_matmul_11_stream_ivalid_2 <= 0;
      __stream_matmul_11_stream_ivalid_3 <= 0;
      __stream_matmul_11_stream_ivalid_4 <= 0;
      __stream_matmul_11_stream_ivalid_5 <= 0;
      __stream_matmul_11_stream_ivalid_6 <= 0;
      __stream_matmul_11_stream_ivalid_7 <= 0;
      __stream_matmul_11_stream_ivalid_8 <= 0;
      __stream_matmul_11_stream_ivalid_9 <= 0;
      __stream_matmul_11_stream_ivalid_10 <= 0;
      __stream_matmul_11_stream_ivalid_11 <= 0;
      __stream_matmul_11_stream_ivalid_12 <= 0;
      __stream_matmul_11_stream_ivalid_13 <= 0;
      __stream_matmul_11_stream_ivalid_14 <= 0;
      __stream_matmul_11_stream_ivalid_15 <= 0;
      __stream_matmul_11_stream_ivalid_16 <= 0;
      __stream_matmul_11_stream_ivalid_17 <= 0;
      __stream_matmul_11_stream_ivalid_18 <= 0;
      __stream_matmul_11_stream_ivalid_19 <= 0;
      __stream_matmul_11_stream_ivalid_20 <= 0;
      __stream_matmul_11_stream_ivalid_21 <= 0;
      __stream_matmul_11_stream_ivalid_22 <= 0;
      __stream_matmul_11_stream_ivalid_23 <= 0;
      __stream_matmul_11_stream_ivalid_24 <= 0;
      __stream_matmul_11_stream_ivalid_25 <= 0;
      __stream_matmul_11_stream_ivalid_26 <= 0;
      __stream_matmul_11_stream_ivalid_27 <= 0;
      __stream_matmul_11_stream_ivalid_28 <= 0;
      __stream_matmul_11_stream_ivalid_29 <= 0;
      _eq_data_2211 <= 0;
      _eq_data_2215 <= 0;
      _plus_data_2235 <= 0;
      _plus_data_2240 <= 0;
      _plus_data_2245 <= 0;
      _eq_data_2251 <= 0;
      _eq_data_2254 <= 0;
      __delay_data_2403__variable_2210 <= 0;
      __delay_data_2404_pointer_2230 <= 0;
      __delay_data_2405_reinterpretcast_2229 <= 0;
      __delay_data_2406__variable_2161 <= 0;
      __delay_data_2427__variable_2156 <= 0;
      __delay_data_2438_cond_2177 <= 0;
      __delay_data_2455_cond_2184 <= 0;
      __delay_data_2407__delay_2406__variable_2161 <= 0;
      __delay_data_2417_plus_2240 <= 0;
      __delay_data_2428__delay_2427__variable_2156 <= 0;
      __delay_data_2439__delay_2438_cond_2177 <= 0;
      __delay_data_2456__delay_2455_cond_2184 <= 0;
      __delay_data_2473_plus_2245 <= 0;
      __delay_data_2491_eq_2251 <= 0;
      __delay_data_2520_eq_2254 <= 0;
      __delay_data_2408__delay_2407__delay_2406__variable_2161 <= 0;
      __delay_data_2418__delay_2417_plus_2240 <= 0;
      __delay_data_2429__delay_2428__delay_2427__variable_2156 <= 0;
      __delay_data_2440__delay_2439__delay_2438_cond_2177 <= 0;
      __delay_data_2457__delay_2456__delay_2455_cond_2184 <= 0;
      __delay_data_2474__delay_2473_plus_2245 <= 0;
      __delay_data_2492__delay_2491_eq_2251 <= 0;
      __delay_data_2521__delay_2520_eq_2254 <= 0;
      __delay_data_2409__delay_2408__delay_2407____variable_2161 <= 0;
      __delay_data_2419__delay_2418__delay_2417_plus_2240 <= 0;
      __delay_data_2430__delay_2429__delay_2428____variable_2156 <= 0;
      __delay_data_2441__delay_2440__delay_2439___cond_2177 <= 0;
      __delay_data_2458__delay_2457__delay_2456___cond_2184 <= 0;
      __delay_data_2475__delay_2474__delay_2473_plus_2245 <= 0;
      __delay_data_2493__delay_2492__delay_2491_eq_2251 <= 0;
      __delay_data_2522__delay_2521__delay_2520_eq_2254 <= 0;
      __delay_data_2410__delay_2409__delay_2408____variable_2161 <= 0;
      __delay_data_2420__delay_2419__delay_2418___plus_2240 <= 0;
      __delay_data_2431__delay_2430__delay_2429____variable_2156 <= 0;
      __delay_data_2442__delay_2441__delay_2440___cond_2177 <= 0;
      __delay_data_2459__delay_2458__delay_2457___cond_2184 <= 0;
      __delay_data_2476__delay_2475__delay_2474___plus_2245 <= 0;
      __delay_data_2494__delay_2493__delay_2492__delay_2491_eq_2251 <= 0;
      __delay_data_2523__delay_2522__delay_2521__delay_2520_eq_2254 <= 0;
      __delay_data_2411__delay_2410__delay_2409____variable_2161 <= 0;
      __delay_data_2421__delay_2420__delay_2419___plus_2240 <= 0;
      __delay_data_2432__delay_2431__delay_2430____variable_2156 <= 0;
      __delay_data_2443__delay_2442__delay_2441___cond_2177 <= 0;
      __delay_data_2460__delay_2459__delay_2458___cond_2184 <= 0;
      __delay_data_2477__delay_2476__delay_2475___plus_2245 <= 0;
      __delay_data_2495__delay_2494__delay_2493__delay_2492___eq_2251 <= 0;
      __delay_data_2524__delay_2523__delay_2522__delay_2521___eq_2254 <= 0;
      __delay_data_2412__delay_2411__delay_2410____variable_2161 <= 0;
      __delay_data_2422__delay_2421__delay_2420___plus_2240 <= 0;
      __delay_data_2433__delay_2432__delay_2431____variable_2156 <= 0;
      __delay_data_2444__delay_2443__delay_2442___cond_2177 <= 0;
      __delay_data_2461__delay_2460__delay_2459___cond_2184 <= 0;
      __delay_data_2478__delay_2477__delay_2476___plus_2245 <= 0;
      __delay_data_2496__delay_2495__delay_2494__delay_2493___eq_2251 <= 0;
      __delay_data_2525__delay_2524__delay_2523__delay_2522___eq_2254 <= 0;
      __delay_data_2413__delay_2412__delay_2411____variable_2161 <= 0;
      __delay_data_2423__delay_2422__delay_2421___plus_2240 <= 0;
      __delay_data_2434__delay_2433__delay_2432____variable_2156 <= 0;
      __delay_data_2445__delay_2444__delay_2443___cond_2177 <= 0;
      __delay_data_2462__delay_2461__delay_2460___cond_2184 <= 0;
      __delay_data_2479__delay_2478__delay_2477___plus_2245 <= 0;
      __delay_data_2497__delay_2496__delay_2495__delay_2494___eq_2251 <= 0;
      __delay_data_2526__delay_2525__delay_2524__delay_2523___eq_2254 <= 0;
      __delay_data_2414__delay_2413__delay_2412____variable_2161 <= 0;
      __delay_data_2424__delay_2423__delay_2422___plus_2240 <= 0;
      __delay_data_2435__delay_2434__delay_2433____variable_2156 <= 0;
      __delay_data_2446__delay_2445__delay_2444___cond_2177 <= 0;
      __delay_data_2463__delay_2462__delay_2461___cond_2184 <= 0;
      __delay_data_2480__delay_2479__delay_2478___plus_2245 <= 0;
      __delay_data_2498__delay_2497__delay_2496__delay_2495___eq_2251 <= 0;
      __delay_data_2527__delay_2526__delay_2525__delay_2524___eq_2254 <= 0;
      __delay_data_2415__delay_2414__delay_2413____variable_2161 <= 0;
      __delay_data_2425__delay_2424__delay_2423___plus_2240 <= 0;
      __delay_data_2436__delay_2435__delay_2434____variable_2156 <= 0;
      __delay_data_2447__delay_2446__delay_2445___cond_2177 <= 0;
      __delay_data_2464__delay_2463__delay_2462___cond_2184 <= 0;
      __delay_data_2481__delay_2480__delay_2479___plus_2245 <= 0;
      __delay_data_2499__delay_2498__delay_2497__delay_2496___eq_2251 <= 0;
      __delay_data_2528__delay_2527__delay_2526__delay_2525___eq_2254 <= 0;
      __delay_data_2416__delay_2415__delay_2414____variable_2161 <= 0;
      __delay_data_2426__delay_2425__delay_2424___plus_2240 <= 0;
      __delay_data_2437__delay_2436__delay_2435____variable_2156 <= 0;
      __delay_data_2448__delay_2447__delay_2446___cond_2177 <= 0;
      __delay_data_2465__delay_2464__delay_2463___cond_2184 <= 0;
      __delay_data_2482__delay_2481__delay_2480___plus_2245 <= 0;
      __delay_data_2500__delay_2499__delay_2498__delay_2497___eq_2251 <= 0;
      __delay_data_2529__delay_2528__delay_2527__delay_2526___eq_2254 <= 0;
      __delay_data_2449__delay_2448__delay_2447___cond_2177 <= 0;
      __delay_data_2466__delay_2465__delay_2464___cond_2184 <= 0;
      __delay_data_2483__delay_2482__delay_2481___plus_2245 <= 0;
      __delay_data_2501__delay_2500__delay_2499__delay_2498___eq_2251 <= 0;
      __delay_data_2530__delay_2529__delay_2528__delay_2527___eq_2254 <= 0;
      __delay_data_2450__delay_2449__delay_2448___cond_2177 <= 0;
      __delay_data_2467__delay_2466__delay_2465___cond_2184 <= 0;
      __delay_data_2484__delay_2483__delay_2482___plus_2245 <= 0;
      __delay_data_2502__delay_2501__delay_2500__delay_2499___eq_2251 <= 0;
      __delay_data_2531__delay_2530__delay_2529__delay_2528___eq_2254 <= 0;
      __delay_data_2451__delay_2450__delay_2449___cond_2177 <= 0;
      __delay_data_2468__delay_2467__delay_2466___cond_2184 <= 0;
      __delay_data_2485__delay_2484__delay_2483___plus_2245 <= 0;
      __delay_data_2503__delay_2502__delay_2501__delay_2500___eq_2251 <= 0;
      __delay_data_2532__delay_2531__delay_2530__delay_2529___eq_2254 <= 0;
      __delay_data_2452__delay_2451__delay_2450___cond_2177 <= 0;
      __delay_data_2469__delay_2468__delay_2467___cond_2184 <= 0;
      __delay_data_2486__delay_2485__delay_2484___plus_2245 <= 0;
      __delay_data_2504__delay_2503__delay_2502__delay_2501___eq_2251 <= 0;
      __delay_data_2533__delay_2532__delay_2531__delay_2530___eq_2254 <= 0;
      __delay_data_2453__delay_2452__delay_2451___cond_2177 <= 0;
      __delay_data_2470__delay_2469__delay_2468___cond_2184 <= 0;
      __delay_data_2487__delay_2486__delay_2485___plus_2245 <= 0;
      __delay_data_2505__delay_2504__delay_2503__delay_2502___eq_2251 <= 0;
      __delay_data_2534__delay_2533__delay_2532__delay_2531___eq_2254 <= 0;
      __delay_data_2454__delay_2453__delay_2452___cond_2177 <= 0;
      __delay_data_2471__delay_2470__delay_2469___cond_2184 <= 0;
      __delay_data_2488__delay_2487__delay_2486___plus_2245 <= 0;
      __delay_data_2506__delay_2505__delay_2504__delay_2503___eq_2251 <= 0;
      __delay_data_2535__delay_2534__delay_2533__delay_2532___eq_2254 <= 0;
      _plus_data_2243 <= 0;
      __delay_data_2472__delay_2471__delay_2470___cond_2184 <= 0;
      __delay_data_2489__delay_2488__delay_2487___plus_2245 <= 0;
      __delay_data_2507__delay_2506__delay_2505__delay_2504___eq_2251 <= 0;
      __delay_data_2536__delay_2535__delay_2534__delay_2533___eq_2254 <= 0;
      __delay_data_2548__substreamoutput_2242 <= 0;
      __delay_data_2508__delay_2507__delay_2506__delay_2505___eq_2251 <= 0;
      __delay_data_2537__delay_2536__delay_2535__delay_2534___eq_2254 <= 0;
      __delay_data_2549__delay_2548__substreamoutput_2242 <= 0;
      __delay_data_2509__delay_2508__delay_2507__delay_2506___eq_2251 <= 0;
      __delay_data_2538__delay_2537__delay_2536__delay_2535___eq_2254 <= 0;
      __delay_data_2550__delay_2549____substreamoutput_2242 <= 0;
      __delay_data_2510__delay_2509__delay_2508__delay_2507___eq_2251 <= 0;
      __delay_data_2539__delay_2538__delay_2537__delay_2536___eq_2254 <= 0;
      __delay_data_2551__delay_2550____substreamoutput_2242 <= 0;
      __delay_data_2511__delay_2510__delay_2509__delay_2508___eq_2251 <= 0;
      __delay_data_2540__delay_2539__delay_2538__delay_2537___eq_2254 <= 0;
      __delay_data_2552__delay_2551____substreamoutput_2242 <= 0;
      __delay_data_2512__delay_2511__delay_2510__delay_2509___eq_2251 <= 0;
      __delay_data_2541__delay_2540__delay_2539__delay_2538___eq_2254 <= 0;
      __delay_data_2553__delay_2552____substreamoutput_2242 <= 0;
      __delay_data_2513__delay_2512__delay_2511__delay_2510___eq_2251 <= 0;
      __delay_data_2542__delay_2541__delay_2540__delay_2539___eq_2254 <= 0;
      __delay_data_2554__delay_2553____substreamoutput_2242 <= 0;
      __delay_data_2514__delay_2513__delay_2512__delay_2511___eq_2251 <= 0;
      __delay_data_2543__delay_2542__delay_2541__delay_2540___eq_2254 <= 0;
      __delay_data_2555__delay_2554____substreamoutput_2242 <= 0;
      __delay_data_2515__delay_2514__delay_2513__delay_2512___eq_2251 <= 0;
      __delay_data_2544__delay_2543__delay_2542__delay_2541___eq_2254 <= 0;
      __delay_data_2556__delay_2555____substreamoutput_2242 <= 0;
      __delay_data_2516__delay_2515__delay_2514__delay_2513___eq_2251 <= 0;
      __delay_data_2545__delay_2544__delay_2543__delay_2542___eq_2254 <= 0;
      __delay_data_2557__delay_2556____substreamoutput_2242 <= 0;
      _greaterthan_data_2248 <= 0;
      __delay_data_2490__substreamoutput_2246 <= 0;
      __delay_data_2517__delay_2516__delay_2515__delay_2514___eq_2251 <= 0;
      __delay_data_2546__delay_2545__delay_2544__delay_2543___eq_2254 <= 0;
      __delay_data_2558__delay_2557____substreamoutput_2242 <= 0;
      _cond_data_2250 <= 0;
      __delay_data_2518__delay_2517__delay_2516__delay_2515___eq_2251 <= 0;
      __delay_data_2519__delay_2490__substreamoutput_2246 <= 0;
      __delay_data_2547__delay_2546__delay_2545__delay_2544___eq_2254 <= 0;
      __delay_data_2559__delay_2558____substreamoutput_2242 <= 0;
      _stream_matmul_11_parameter_0_next_parameter_data <= 0;
      __variable_wdata_2156 <= 0;
      _stream_matmul_11_parameter_1_next_parameter_data <= 0;
      __variable_wdata_2157 <= 0;
      _stream_matmul_11_parameter_2_next_parameter_data <= 0;
      __variable_wdata_2158 <= 0;
      _stream_matmul_11_parameter_3_next_parameter_data <= 0;
      __variable_wdata_2159 <= 0;
      _stream_matmul_11_parameter_4_next_parameter_data <= 0;
      __variable_wdata_2160 <= 0;
      _stream_matmul_11_parameter_6_next_parameter_data <= 0;
      __variable_wdata_2171 <= 0;
      _stream_matmul_11_source_7_source_mode <= 5'b0;
      _stream_matmul_11_source_7_source_offset <= 0;
      _source_stream_matmul_11_source_7_pat_size_0 <= 0;
      _source_stream_matmul_11_source_7_pat_stride_0 <= 0;
      _source_stream_matmul_11_source_7_pat_size_1 <= 0;
      _source_stream_matmul_11_source_7_pat_stride_1 <= 0;
      _source_stream_matmul_11_source_7_pat_size_2 <= 0;
      _source_stream_matmul_11_source_7_pat_stride_2 <= 0;
      _source_stream_matmul_11_source_7_pat_size_3 <= 0;
      _source_stream_matmul_11_source_7_pat_stride_3 <= 0;
      _stream_matmul_11_source_7_source_sel <= 0;
      _stream_matmul_11_source_7_source_offset_buf <= 0;
      _source_stream_matmul_11_source_7_pat_cur_offset_0 <= 0;
      _source_stream_matmul_11_source_7_pat_cur_offset_1 <= 0;
      _source_stream_matmul_11_source_7_pat_cur_offset_2 <= 0;
      _source_stream_matmul_11_source_7_pat_cur_offset_3 <= 0;
      _source_stream_matmul_11_source_7_pat_count_0 <= 0;
      _source_stream_matmul_11_source_7_pat_count_1 <= 0;
      _source_stream_matmul_11_source_7_pat_count_2 <= 0;
      _source_stream_matmul_11_source_7_pat_count_3 <= 0;
      _source_stream_matmul_11_source_7_pat_size_buf_0 <= 0;
      _source_stream_matmul_11_source_7_pat_size_buf_1 <= 0;
      _source_stream_matmul_11_source_7_pat_size_buf_2 <= 0;
      _source_stream_matmul_11_source_7_pat_size_buf_3 <= 0;
      _source_stream_matmul_11_source_7_pat_stride_buf_0 <= 0;
      _source_stream_matmul_11_source_7_pat_stride_buf_1 <= 0;
      _source_stream_matmul_11_source_7_pat_stride_buf_2 <= 0;
      _source_stream_matmul_11_source_7_pat_stride_buf_3 <= 0;
      __variable_wdata_2172 <= 0;
      _stream_matmul_11_source_7_source_ram_raddr <= 0;
      _stream_matmul_11_parameter_8_next_parameter_data <= 0;
      __variable_wdata_2178 <= 0;
      _stream_matmul_11_source_9_source_mode <= 5'b0;
      _stream_matmul_11_source_9_source_offset <= 0;
      _source_stream_matmul_11_source_9_pat_size_0 <= 0;
      _source_stream_matmul_11_source_9_pat_stride_0 <= 0;
      _source_stream_matmul_11_source_9_pat_size_1 <= 0;
      _source_stream_matmul_11_source_9_pat_stride_1 <= 0;
      _source_stream_matmul_11_source_9_pat_size_2 <= 0;
      _source_stream_matmul_11_source_9_pat_stride_2 <= 0;
      _source_stream_matmul_11_source_9_pat_size_3 <= 0;
      _source_stream_matmul_11_source_9_pat_stride_3 <= 0;
      _stream_matmul_11_source_9_source_sel <= 0;
      _stream_matmul_11_source_9_source_offset_buf <= 0;
      _source_stream_matmul_11_source_9_pat_cur_offset_0 <= 0;
      _source_stream_matmul_11_source_9_pat_cur_offset_1 <= 0;
      _source_stream_matmul_11_source_9_pat_cur_offset_2 <= 0;
      _source_stream_matmul_11_source_9_pat_cur_offset_3 <= 0;
      _source_stream_matmul_11_source_9_pat_count_0 <= 0;
      _source_stream_matmul_11_source_9_pat_count_1 <= 0;
      _source_stream_matmul_11_source_9_pat_count_2 <= 0;
      _source_stream_matmul_11_source_9_pat_count_3 <= 0;
      _source_stream_matmul_11_source_9_pat_size_buf_0 <= 0;
      _source_stream_matmul_11_source_9_pat_size_buf_1 <= 0;
      _source_stream_matmul_11_source_9_pat_size_buf_2 <= 0;
      _source_stream_matmul_11_source_9_pat_size_buf_3 <= 0;
      _source_stream_matmul_11_source_9_pat_stride_buf_0 <= 0;
      _source_stream_matmul_11_source_9_pat_stride_buf_1 <= 0;
      _source_stream_matmul_11_source_9_pat_stride_buf_2 <= 0;
      _source_stream_matmul_11_source_9_pat_stride_buf_3 <= 0;
      __variable_wdata_2179 <= 0;
      _stream_matmul_11_source_9_source_ram_raddr <= 0;
      _stream_matmul_11_parameter_10_next_parameter_data <= 0;
      __variable_wdata_2185 <= 0;
      _stream_matmul_11_source_11_source_mode <= 5'b0;
      _stream_matmul_11_source_11_source_empty_data <= 0;
      __variable_wdata_2186 <= 0;
      _stream_matmul_11_parameter_12_next_parameter_data <= 0;
      __variable_wdata_2192 <= 0;
      _stream_matmul_11_source_13_source_mode <= 5'b0;
      _stream_matmul_11_source_13_source_empty_data <= 0;
      __variable_wdata_2193 <= 0;
      _stream_matmul_11_parameter_14_next_parameter_data <= 0;
      __variable_wdata_2199 <= 0;
      _stream_matmul_11_source_15_source_mode <= 5'b0;
      _stream_matmul_11_source_15_source_empty_data <= 0;
      __variable_wdata_2200 <= 0;
      _stream_matmul_11_parameter_16_next_parameter_data <= 0;
      __variable_wdata_2206 <= 0;
      _stream_matmul_11_parameter_17_next_parameter_data <= 0;
      __variable_wdata_2207 <= 0;
      _stream_matmul_11_parameter_18_next_parameter_data <= 0;
      __variable_wdata_2208 <= 0;
      _stream_matmul_11_parameter_19_next_parameter_data <= 0;
      __variable_wdata_2209 <= 0;
      _stream_matmul_11_source_20_source_mode <= 5'b0;
      _stream_matmul_11_source_20_source_offset <= 0;
      _source_stream_matmul_11_source_20_pat_size_0 <= 0;
      _source_stream_matmul_11_source_20_pat_stride_0 <= 0;
      _source_stream_matmul_11_source_20_pat_size_1 <= 0;
      _source_stream_matmul_11_source_20_pat_stride_1 <= 0;
      _source_stream_matmul_11_source_20_pat_size_2 <= 0;
      _source_stream_matmul_11_source_20_pat_stride_2 <= 0;
      _source_stream_matmul_11_source_20_pat_size_3 <= 0;
      _source_stream_matmul_11_source_20_pat_stride_3 <= 0;
      _stream_matmul_11_source_20_source_sel <= 0;
      _stream_matmul_11_source_20_source_offset_buf <= 0;
      _source_stream_matmul_11_source_20_pat_cur_offset_0 <= 0;
      _source_stream_matmul_11_source_20_pat_cur_offset_1 <= 0;
      _source_stream_matmul_11_source_20_pat_cur_offset_2 <= 0;
      _source_stream_matmul_11_source_20_pat_cur_offset_3 <= 0;
      _source_stream_matmul_11_source_20_pat_count_0 <= 0;
      _source_stream_matmul_11_source_20_pat_count_1 <= 0;
      _source_stream_matmul_11_source_20_pat_count_2 <= 0;
      _source_stream_matmul_11_source_20_pat_count_3 <= 0;
      _source_stream_matmul_11_source_20_pat_size_buf_0 <= 0;
      _source_stream_matmul_11_source_20_pat_size_buf_1 <= 0;
      _source_stream_matmul_11_source_20_pat_size_buf_2 <= 0;
      _source_stream_matmul_11_source_20_pat_size_buf_3 <= 0;
      _source_stream_matmul_11_source_20_pat_stride_buf_0 <= 0;
      _source_stream_matmul_11_source_20_pat_stride_buf_1 <= 0;
      _source_stream_matmul_11_source_20_pat_stride_buf_2 <= 0;
      _source_stream_matmul_11_source_20_pat_stride_buf_3 <= 0;
      __variable_wdata_2210 <= 0;
      _stream_matmul_11_source_20_source_ram_raddr <= 0;
      _stream_matmul_11_source_21_source_mode <= 5'b0;
      _stream_matmul_11_source_21_source_offset <= 0;
      _source_stream_matmul_11_source_21_pat_size_0 <= 0;
      _source_stream_matmul_11_source_21_pat_stride_0 <= 0;
      _source_stream_matmul_11_source_21_pat_size_1 <= 0;
      _source_stream_matmul_11_source_21_pat_stride_1 <= 0;
      _source_stream_matmul_11_source_21_pat_size_2 <= 0;
      _source_stream_matmul_11_source_21_pat_stride_2 <= 0;
      _source_stream_matmul_11_source_21_pat_size_3 <= 0;
      _source_stream_matmul_11_source_21_pat_stride_3 <= 0;
      _stream_matmul_11_source_21_source_sel <= 0;
      _stream_matmul_11_source_21_source_offset_buf <= 0;
      _source_stream_matmul_11_source_21_pat_cur_offset_0 <= 0;
      _source_stream_matmul_11_source_21_pat_cur_offset_1 <= 0;
      _source_stream_matmul_11_source_21_pat_cur_offset_2 <= 0;
      _source_stream_matmul_11_source_21_pat_cur_offset_3 <= 0;
      _source_stream_matmul_11_source_21_pat_count_0 <= 0;
      _source_stream_matmul_11_source_21_pat_count_1 <= 0;
      _source_stream_matmul_11_source_21_pat_count_2 <= 0;
      _source_stream_matmul_11_source_21_pat_count_3 <= 0;
      _source_stream_matmul_11_source_21_pat_size_buf_0 <= 0;
      _source_stream_matmul_11_source_21_pat_size_buf_1 <= 0;
      _source_stream_matmul_11_source_21_pat_size_buf_2 <= 0;
      _source_stream_matmul_11_source_21_pat_size_buf_3 <= 0;
      _source_stream_matmul_11_source_21_pat_stride_buf_0 <= 0;
      _source_stream_matmul_11_source_21_pat_stride_buf_1 <= 0;
      _source_stream_matmul_11_source_21_pat_stride_buf_2 <= 0;
      _source_stream_matmul_11_source_21_pat_stride_buf_3 <= 0;
      __variable_wdata_2224 <= 0;
      _stream_matmul_11_source_21_source_ram_raddr <= 0;
      _tmp_1410 <= 0;
      _tmp_1411 <= 0;
      _tmp_1412 <= 0;
      _tmp_1413 <= 0;
      _tmp_1414 <= 0;
      _tmp_1415 <= 0;
      _tmp_1416 <= 0;
      _tmp_1417 <= 0;
      _tmp_1418 <= 0;
      _tmp_1419 <= 0;
      _tmp_1420 <= 0;
      _tmp_1421 <= 0;
      _tmp_1422 <= 0;
      _tmp_1423 <= 0;
      _tmp_1424 <= 0;
      _tmp_1425 <= 0;
      _tmp_1426 <= 0;
      _tmp_1427 <= 0;
      _tmp_1428 <= 0;
      _tmp_1429 <= 0;
      _tmp_1430 <= 0;
      _tmp_1431 <= 0;
      _tmp_1432 <= 0;
      _tmp_1433 <= 0;
      _tmp_1434 <= 0;
      _tmp_1435 <= 0;
      _tmp_1436 <= 0;
      _tmp_1437 <= 0;
      _tmp_1438 <= 0;
      _tmp_1439 <= 0;
      _tmp_1440 <= 0;
      _tmp_1443 <= 0;
      _tmp_1444 <= 0;
      _tmp_1445 <= 0;
      _tmp_1446 <= 0;
      _tmp_1447 <= 0;
      _tmp_1448 <= 0;
      _tmp_1449 <= 0;
      _tmp_1450 <= 0;
      _tmp_1451 <= 0;
      _tmp_1452 <= 0;
      _tmp_1453 <= 0;
      _tmp_1454 <= 0;
      _tmp_1455 <= 0;
      _tmp_1456 <= 0;
      _tmp_1457 <= 0;
      _tmp_1458 <= 0;
      _tmp_1459 <= 0;
      _tmp_1460 <= 0;
      _tmp_1461 <= 0;
      _tmp_1462 <= 0;
      _tmp_1463 <= 0;
      _tmp_1464 <= 0;
      _tmp_1465 <= 0;
      _tmp_1466 <= 0;
      _tmp_1467 <= 0;
      _tmp_1468 <= 0;
      _tmp_1469 <= 0;
      _tmp_1470 <= 0;
      _tmp_1471 <= 0;
      _tmp_1472 <= 0;
      _tmp_1473 <= 0;
      _tmp_1474 <= 0;
      _tmp_1475 <= 0;
      _tmp_1476 <= 0;
      _tmp_1477 <= 0;
      _tmp_1478 <= 0;
      _tmp_1479 <= 0;
      _tmp_1480 <= 0;
      _tmp_1481 <= 0;
      _tmp_1482 <= 0;
      _tmp_1483 <= 0;
      _tmp_1484 <= 0;
      _tmp_1485 <= 0;
      _tmp_1486 <= 0;
      _tmp_1487 <= 0;
      _tmp_1488 <= 0;
      _tmp_1489 <= 0;
      _tmp_1490 <= 0;
      _tmp_1491 <= 0;
      _tmp_1492 <= 0;
      _tmp_1493 <= 0;
      _tmp_1494 <= 0;
      _tmp_1495 <= 0;
      _tmp_1496 <= 0;
      _tmp_1497 <= 0;
      _tmp_1498 <= 0;
      _tmp_1499 <= 0;
      _tmp_1500 <= 0;
      _tmp_1501 <= 0;
      _tmp_1502 <= 0;
      _tmp_1503 <= 0;
      _tmp_1504 <= 0;
      _stream_matmul_11_sink_26_sink_mode <= 5'b0;
      _stream_matmul_11_sink_26_sink_offset <= 0;
      _stream_matmul_11_sink_26_sink_size <= 0;
      _stream_matmul_11_sink_26_sink_stride <= 0;
      _stream_matmul_11_sink_26_sink_sel <= 0;
      _stream_matmul_11_sink_26_sink_offset_buf <= 0;
      _stream_matmul_11_sink_26_sink_size_buf <= 0;
      _stream_matmul_11_sink_26_sink_stride_buf <= 0;
      _stream_matmul_11_sink_26_sink_waddr <= 0;
      _stream_matmul_11_sink_26_sink_count <= 0;
      _stream_matmul_11_sink_26_sink_wdata <= 0;
      _tmp_1517 <= 0;
      _tmp_1518 <= 0;
      _tmp_1519 <= 0;
      _tmp_1520 <= 0;
      _tmp_1521 <= 0;
      _tmp_1522 <= 0;
      __variable_wdata_2161 <= 0;
      _tmp_1523 <= 0;
      _tmp_1524 <= 0;
      _tmp_1525 <= 0;
      _tmp_1526 <= 0;
      _tmp_1529 <= 0;
      _tmp_1532 <= 0;
      _tmp_1533 <= 0;
      _tmp_1534 <= 0;
      _tmp_1535 <= 0;
      _tmp_1536 <= 0;
      _tmp_1537 <= 0;
      _tmp_1538 <= 0;
      _tmp_1539 <= 0;
      _tmp_1540 <= 0;
      _tmp_1541 <= 0;
      _tmp_1542 <= 0;
      _tmp_1543 <= 0;
      _tmp_1544 <= 0;
      _tmp_1545 <= 0;
      _tmp_1546 <= 0;
      _tmp_1547 <= 0;
      _tmp_1548 <= 0;
      _tmp_1549 <= 0;
      _tmp_1550 <= 0;
      _tmp_1551 <= 0;
      _tmp_1552 <= 0;
      _tmp_1553 <= 0;
      _tmp_1554 <= 0;
      _tmp_1555 <= 0;
      _tmp_1556 <= 0;
      _tmp_1557 <= 0;
      _tmp_1558 <= 0;
      _tmp_1559 <= 0;
      _tmp_1560 <= 0;
      _tmp_1561 <= 0;
      _tmp_1562 <= 0;
      _tmp_1563 <= 0;
      _tmp_1564 <= 0;
      _tmp_1565 <= 0;
      _tmp_1566 <= 0;
      _tmp_1567 <= 0;
      _tmp_1568 <= 0;
      _tmp_1569 <= 0;
      _tmp_1570 <= 0;
      _tmp_1571 <= 0;
      _tmp_1572 <= 0;
      _tmp_1573 <= 0;
      _tmp_1574 <= 0;
      _tmp_1575 <= 0;
      _tmp_1576 <= 0;
      _tmp_1577 <= 0;
      _tmp_1578 <= 0;
      _tmp_1579 <= 0;
      _tmp_1580 <= 0;
      _tmp_1581 <= 0;
      _tmp_1582 <= 0;
      _tmp_1583 <= 0;
      _tmp_1584 <= 0;
      _tmp_1585 <= 0;
      _tmp_1586 <= 0;
      _tmp_1587 <= 0;
      _tmp_1588 <= 0;
      _tmp_1589 <= 0;
      _tmp_1590 <= 0;
      _tmp_1591 <= 0;
      _tmp_1592 <= 0;
      _tmp_1593 <= 0;
      _tmp_1594 <= 0;
      _tmp_1595 <= 0;
      _tmp_1596 <= 0;
      _tmp_1597 <= 0;
      _tmp_1598 <= 0;
      _tmp_1599 <= 0;
      _tmp_1600 <= 0;
      _tmp_1601 <= 0;
      _tmp_1602 <= 0;
      _tmp_1603 <= 0;
      _tmp_1604 <= 0;
      _tmp_1605 <= 0;
      _tmp_1606 <= 0;
      _tmp_1607 <= 0;
      _tmp_1608 <= 0;
      _tmp_1609 <= 0;
      _tmp_1610 <= 0;
      _tmp_1611 <= 0;
      _tmp_1612 <= 0;
      _tmp_1613 <= 0;
      _tmp_1614 <= 0;
      _tmp_1615 <= 0;
      _tmp_1616 <= 0;
      _tmp_1617 <= 0;
      _tmp_1618 <= 0;
      _tmp_1619 <= 0;
      _tmp_1620 <= 0;
      _tmp_1621 <= 0;
      _tmp_1622 <= 0;
      _tmp_1623 <= 0;
      _tmp_1624 <= 0;
      _tmp_1625 <= 0;
      _tmp_1626 <= 0;
      _stream_matmul_11_busy_reg <= 0;
    end else begin
      if(_stream_matmul_11_stream_oready) begin
        _stream_matmul_11_source_7_source_ram_renable <= 0;
        _stream_matmul_11_source_7_source_fifo_deq <= 0;
      end 
      _stream_matmul_11_source_7_idle <= _stream_matmul_11_source_7_idle;
      if(_stream_matmul_11_stream_oready) begin
        _stream_matmul_11_source_9_source_ram_renable <= 0;
        _stream_matmul_11_source_9_source_fifo_deq <= 0;
      end 
      _stream_matmul_11_source_9_idle <= _stream_matmul_11_source_9_idle;
      if(_stream_matmul_11_stream_oready) begin
        _stream_matmul_11_source_11_source_ram_renable <= 0;
        _stream_matmul_11_source_11_source_fifo_deq <= 0;
      end 
      _stream_matmul_11_source_11_idle <= _stream_matmul_11_source_11_idle;
      if(_stream_matmul_11_stream_oready) begin
        _stream_matmul_11_source_13_source_ram_renable <= 0;
        _stream_matmul_11_source_13_source_fifo_deq <= 0;
      end 
      _stream_matmul_11_source_13_idle <= _stream_matmul_11_source_13_idle;
      if(_stream_matmul_11_stream_oready) begin
        _stream_matmul_11_source_15_source_ram_renable <= 0;
        _stream_matmul_11_source_15_source_fifo_deq <= 0;
      end 
      _stream_matmul_11_source_15_idle <= _stream_matmul_11_source_15_idle;
      if(_stream_matmul_11_stream_oready) begin
        _stream_matmul_11_source_20_source_ram_renable <= 0;
        _stream_matmul_11_source_20_source_fifo_deq <= 0;
      end 
      _stream_matmul_11_source_20_idle <= _stream_matmul_11_source_20_idle;
      if(_stream_matmul_11_stream_oready) begin
        _stream_matmul_11_source_21_source_ram_renable <= 0;
        _stream_matmul_11_source_21_source_fifo_deq <= 0;
      end 
      _stream_matmul_11_source_21_idle <= _stream_matmul_11_source_21_idle;
      if(_stream_matmul_11_stream_oready) begin
        _stream_matmul_11_sink_26_sink_wenable <= 0;
        _stream_matmul_11_sink_26_sink_fifo_enq <= 0;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _stream_matmul_11_sink_27_sink_wenable <= 0;
        _stream_matmul_11_sink_27_sink_fifo_enq <= 0;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __stream_matmul_11_stream_ivalid_1 <= _stream_matmul_11_stream_ivalid;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __stream_matmul_11_stream_ivalid_2 <= __stream_matmul_11_stream_ivalid_1;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __stream_matmul_11_stream_ivalid_3 <= __stream_matmul_11_stream_ivalid_2;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __stream_matmul_11_stream_ivalid_4 <= __stream_matmul_11_stream_ivalid_3;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __stream_matmul_11_stream_ivalid_5 <= __stream_matmul_11_stream_ivalid_4;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __stream_matmul_11_stream_ivalid_6 <= __stream_matmul_11_stream_ivalid_5;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __stream_matmul_11_stream_ivalid_7 <= __stream_matmul_11_stream_ivalid_6;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __stream_matmul_11_stream_ivalid_8 <= __stream_matmul_11_stream_ivalid_7;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __stream_matmul_11_stream_ivalid_9 <= __stream_matmul_11_stream_ivalid_8;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __stream_matmul_11_stream_ivalid_10 <= __stream_matmul_11_stream_ivalid_9;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __stream_matmul_11_stream_ivalid_11 <= __stream_matmul_11_stream_ivalid_10;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __stream_matmul_11_stream_ivalid_12 <= __stream_matmul_11_stream_ivalid_11;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __stream_matmul_11_stream_ivalid_13 <= __stream_matmul_11_stream_ivalid_12;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __stream_matmul_11_stream_ivalid_14 <= __stream_matmul_11_stream_ivalid_13;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __stream_matmul_11_stream_ivalid_15 <= __stream_matmul_11_stream_ivalid_14;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __stream_matmul_11_stream_ivalid_16 <= __stream_matmul_11_stream_ivalid_15;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __stream_matmul_11_stream_ivalid_17 <= __stream_matmul_11_stream_ivalid_16;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __stream_matmul_11_stream_ivalid_18 <= __stream_matmul_11_stream_ivalid_17;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __stream_matmul_11_stream_ivalid_19 <= __stream_matmul_11_stream_ivalid_18;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __stream_matmul_11_stream_ivalid_20 <= __stream_matmul_11_stream_ivalid_19;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __stream_matmul_11_stream_ivalid_21 <= __stream_matmul_11_stream_ivalid_20;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __stream_matmul_11_stream_ivalid_22 <= __stream_matmul_11_stream_ivalid_21;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __stream_matmul_11_stream_ivalid_23 <= __stream_matmul_11_stream_ivalid_22;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __stream_matmul_11_stream_ivalid_24 <= __stream_matmul_11_stream_ivalid_23;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __stream_matmul_11_stream_ivalid_25 <= __stream_matmul_11_stream_ivalid_24;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __stream_matmul_11_stream_ivalid_26 <= __stream_matmul_11_stream_ivalid_25;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __stream_matmul_11_stream_ivalid_27 <= __stream_matmul_11_stream_ivalid_26;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __stream_matmul_11_stream_ivalid_28 <= __stream_matmul_11_stream_ivalid_27;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __stream_matmul_11_stream_ivalid_29 <= __stream_matmul_11_stream_ivalid_28;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _eq_data_2211 <= stream_matmul_11_parameter_1_data == 1'sd0;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _eq_data_2215 <= stream_matmul_11_parameter_2_data == 1'sd0;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _plus_data_2235 <= _cond_data_2191 + stream_matmul_11_parameter_16_data;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _plus_data_2240 <= _cond_data_2198 + stream_matmul_11_parameter_17_data;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _plus_data_2245 <= _cond_data_2205 + stream_matmul_11_parameter_18_data;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _eq_data_2251 <= stream_matmul_11_parameter_19_data == 1'sd0;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _eq_data_2254 <= stream_matmul_11_parameter_19_data == 2'sd1;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2403__variable_2210 <= stream_matmul_11_source_20_data;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2404_pointer_2230 <= _pointer_data_2230;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2405_reinterpretcast_2229 <= _reinterpretcast_data_2229;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2406__variable_2161 <= stream_matmul_11__reduce_reset_data;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2427__variable_2156 <= stream_matmul_11_parameter_0_data;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2438_cond_2177 <= _cond_data_2177;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2455_cond_2184 <= _cond_data_2184;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2407__delay_2406__variable_2161 <= __delay_data_2406__variable_2161;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2417_plus_2240 <= _plus_data_2240;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2428__delay_2427__variable_2156 <= __delay_data_2427__variable_2156;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2439__delay_2438_cond_2177 <= __delay_data_2438_cond_2177;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2456__delay_2455_cond_2184 <= __delay_data_2455_cond_2184;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2473_plus_2245 <= _plus_data_2245;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2491_eq_2251 <= _eq_data_2251;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2520_eq_2254 <= _eq_data_2254;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2408__delay_2407__delay_2406__variable_2161 <= __delay_data_2407__delay_2406__variable_2161;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2418__delay_2417_plus_2240 <= __delay_data_2417_plus_2240;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2429__delay_2428__delay_2427__variable_2156 <= __delay_data_2428__delay_2427__variable_2156;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2440__delay_2439__delay_2438_cond_2177 <= __delay_data_2439__delay_2438_cond_2177;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2457__delay_2456__delay_2455_cond_2184 <= __delay_data_2456__delay_2455_cond_2184;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2474__delay_2473_plus_2245 <= __delay_data_2473_plus_2245;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2492__delay_2491_eq_2251 <= __delay_data_2491_eq_2251;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2521__delay_2520_eq_2254 <= __delay_data_2520_eq_2254;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2409__delay_2408__delay_2407____variable_2161 <= __delay_data_2408__delay_2407__delay_2406__variable_2161;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2419__delay_2418__delay_2417_plus_2240 <= __delay_data_2418__delay_2417_plus_2240;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2430__delay_2429__delay_2428____variable_2156 <= __delay_data_2429__delay_2428__delay_2427__variable_2156;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2441__delay_2440__delay_2439___cond_2177 <= __delay_data_2440__delay_2439__delay_2438_cond_2177;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2458__delay_2457__delay_2456___cond_2184 <= __delay_data_2457__delay_2456__delay_2455_cond_2184;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2475__delay_2474__delay_2473_plus_2245 <= __delay_data_2474__delay_2473_plus_2245;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2493__delay_2492__delay_2491_eq_2251 <= __delay_data_2492__delay_2491_eq_2251;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2522__delay_2521__delay_2520_eq_2254 <= __delay_data_2521__delay_2520_eq_2254;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2410__delay_2409__delay_2408____variable_2161 <= __delay_data_2409__delay_2408__delay_2407____variable_2161;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2420__delay_2419__delay_2418___plus_2240 <= __delay_data_2419__delay_2418__delay_2417_plus_2240;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2431__delay_2430__delay_2429____variable_2156 <= __delay_data_2430__delay_2429__delay_2428____variable_2156;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2442__delay_2441__delay_2440___cond_2177 <= __delay_data_2441__delay_2440__delay_2439___cond_2177;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2459__delay_2458__delay_2457___cond_2184 <= __delay_data_2458__delay_2457__delay_2456___cond_2184;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2476__delay_2475__delay_2474___plus_2245 <= __delay_data_2475__delay_2474__delay_2473_plus_2245;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2494__delay_2493__delay_2492__delay_2491_eq_2251 <= __delay_data_2493__delay_2492__delay_2491_eq_2251;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2523__delay_2522__delay_2521__delay_2520_eq_2254 <= __delay_data_2522__delay_2521__delay_2520_eq_2254;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2411__delay_2410__delay_2409____variable_2161 <= __delay_data_2410__delay_2409__delay_2408____variable_2161;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2421__delay_2420__delay_2419___plus_2240 <= __delay_data_2420__delay_2419__delay_2418___plus_2240;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2432__delay_2431__delay_2430____variable_2156 <= __delay_data_2431__delay_2430__delay_2429____variable_2156;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2443__delay_2442__delay_2441___cond_2177 <= __delay_data_2442__delay_2441__delay_2440___cond_2177;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2460__delay_2459__delay_2458___cond_2184 <= __delay_data_2459__delay_2458__delay_2457___cond_2184;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2477__delay_2476__delay_2475___plus_2245 <= __delay_data_2476__delay_2475__delay_2474___plus_2245;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2495__delay_2494__delay_2493__delay_2492___eq_2251 <= __delay_data_2494__delay_2493__delay_2492__delay_2491_eq_2251;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2524__delay_2523__delay_2522__delay_2521___eq_2254 <= __delay_data_2523__delay_2522__delay_2521__delay_2520_eq_2254;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2412__delay_2411__delay_2410____variable_2161 <= __delay_data_2411__delay_2410__delay_2409____variable_2161;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2422__delay_2421__delay_2420___plus_2240 <= __delay_data_2421__delay_2420__delay_2419___plus_2240;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2433__delay_2432__delay_2431____variable_2156 <= __delay_data_2432__delay_2431__delay_2430____variable_2156;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2444__delay_2443__delay_2442___cond_2177 <= __delay_data_2443__delay_2442__delay_2441___cond_2177;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2461__delay_2460__delay_2459___cond_2184 <= __delay_data_2460__delay_2459__delay_2458___cond_2184;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2478__delay_2477__delay_2476___plus_2245 <= __delay_data_2477__delay_2476__delay_2475___plus_2245;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2496__delay_2495__delay_2494__delay_2493___eq_2251 <= __delay_data_2495__delay_2494__delay_2493__delay_2492___eq_2251;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2525__delay_2524__delay_2523__delay_2522___eq_2254 <= __delay_data_2524__delay_2523__delay_2522__delay_2521___eq_2254;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2413__delay_2412__delay_2411____variable_2161 <= __delay_data_2412__delay_2411__delay_2410____variable_2161;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2423__delay_2422__delay_2421___plus_2240 <= __delay_data_2422__delay_2421__delay_2420___plus_2240;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2434__delay_2433__delay_2432____variable_2156 <= __delay_data_2433__delay_2432__delay_2431____variable_2156;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2445__delay_2444__delay_2443___cond_2177 <= __delay_data_2444__delay_2443__delay_2442___cond_2177;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2462__delay_2461__delay_2460___cond_2184 <= __delay_data_2461__delay_2460__delay_2459___cond_2184;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2479__delay_2478__delay_2477___plus_2245 <= __delay_data_2478__delay_2477__delay_2476___plus_2245;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2497__delay_2496__delay_2495__delay_2494___eq_2251 <= __delay_data_2496__delay_2495__delay_2494__delay_2493___eq_2251;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2526__delay_2525__delay_2524__delay_2523___eq_2254 <= __delay_data_2525__delay_2524__delay_2523__delay_2522___eq_2254;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2414__delay_2413__delay_2412____variable_2161 <= __delay_data_2413__delay_2412__delay_2411____variable_2161;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2424__delay_2423__delay_2422___plus_2240 <= __delay_data_2423__delay_2422__delay_2421___plus_2240;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2435__delay_2434__delay_2433____variable_2156 <= __delay_data_2434__delay_2433__delay_2432____variable_2156;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2446__delay_2445__delay_2444___cond_2177 <= __delay_data_2445__delay_2444__delay_2443___cond_2177;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2463__delay_2462__delay_2461___cond_2184 <= __delay_data_2462__delay_2461__delay_2460___cond_2184;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2480__delay_2479__delay_2478___plus_2245 <= __delay_data_2479__delay_2478__delay_2477___plus_2245;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2498__delay_2497__delay_2496__delay_2495___eq_2251 <= __delay_data_2497__delay_2496__delay_2495__delay_2494___eq_2251;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2527__delay_2526__delay_2525__delay_2524___eq_2254 <= __delay_data_2526__delay_2525__delay_2524__delay_2523___eq_2254;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2415__delay_2414__delay_2413____variable_2161 <= __delay_data_2414__delay_2413__delay_2412____variable_2161;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2425__delay_2424__delay_2423___plus_2240 <= __delay_data_2424__delay_2423__delay_2422___plus_2240;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2436__delay_2435__delay_2434____variable_2156 <= __delay_data_2435__delay_2434__delay_2433____variable_2156;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2447__delay_2446__delay_2445___cond_2177 <= __delay_data_2446__delay_2445__delay_2444___cond_2177;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2464__delay_2463__delay_2462___cond_2184 <= __delay_data_2463__delay_2462__delay_2461___cond_2184;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2481__delay_2480__delay_2479___plus_2245 <= __delay_data_2480__delay_2479__delay_2478___plus_2245;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2499__delay_2498__delay_2497__delay_2496___eq_2251 <= __delay_data_2498__delay_2497__delay_2496__delay_2495___eq_2251;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2528__delay_2527__delay_2526__delay_2525___eq_2254 <= __delay_data_2527__delay_2526__delay_2525__delay_2524___eq_2254;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2416__delay_2415__delay_2414____variable_2161 <= __delay_data_2415__delay_2414__delay_2413____variable_2161;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2426__delay_2425__delay_2424___plus_2240 <= __delay_data_2425__delay_2424__delay_2423___plus_2240;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2437__delay_2436__delay_2435____variable_2156 <= __delay_data_2436__delay_2435__delay_2434____variable_2156;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2448__delay_2447__delay_2446___cond_2177 <= __delay_data_2447__delay_2446__delay_2445___cond_2177;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2465__delay_2464__delay_2463___cond_2184 <= __delay_data_2464__delay_2463__delay_2462___cond_2184;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2482__delay_2481__delay_2480___plus_2245 <= __delay_data_2481__delay_2480__delay_2479___plus_2245;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2500__delay_2499__delay_2498__delay_2497___eq_2251 <= __delay_data_2499__delay_2498__delay_2497__delay_2496___eq_2251;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2529__delay_2528__delay_2527__delay_2526___eq_2254 <= __delay_data_2528__delay_2527__delay_2526__delay_2525___eq_2254;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2449__delay_2448__delay_2447___cond_2177 <= __delay_data_2448__delay_2447__delay_2446___cond_2177;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2466__delay_2465__delay_2464___cond_2184 <= __delay_data_2465__delay_2464__delay_2463___cond_2184;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2483__delay_2482__delay_2481___plus_2245 <= __delay_data_2482__delay_2481__delay_2480___plus_2245;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2501__delay_2500__delay_2499__delay_2498___eq_2251 <= __delay_data_2500__delay_2499__delay_2498__delay_2497___eq_2251;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2530__delay_2529__delay_2528__delay_2527___eq_2254 <= __delay_data_2529__delay_2528__delay_2527__delay_2526___eq_2254;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2450__delay_2449__delay_2448___cond_2177 <= __delay_data_2449__delay_2448__delay_2447___cond_2177;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2467__delay_2466__delay_2465___cond_2184 <= __delay_data_2466__delay_2465__delay_2464___cond_2184;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2484__delay_2483__delay_2482___plus_2245 <= __delay_data_2483__delay_2482__delay_2481___plus_2245;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2502__delay_2501__delay_2500__delay_2499___eq_2251 <= __delay_data_2501__delay_2500__delay_2499__delay_2498___eq_2251;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2531__delay_2530__delay_2529__delay_2528___eq_2254 <= __delay_data_2530__delay_2529__delay_2528__delay_2527___eq_2254;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2451__delay_2450__delay_2449___cond_2177 <= __delay_data_2450__delay_2449__delay_2448___cond_2177;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2468__delay_2467__delay_2466___cond_2184 <= __delay_data_2467__delay_2466__delay_2465___cond_2184;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2485__delay_2484__delay_2483___plus_2245 <= __delay_data_2484__delay_2483__delay_2482___plus_2245;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2503__delay_2502__delay_2501__delay_2500___eq_2251 <= __delay_data_2502__delay_2501__delay_2500__delay_2499___eq_2251;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2532__delay_2531__delay_2530__delay_2529___eq_2254 <= __delay_data_2531__delay_2530__delay_2529__delay_2528___eq_2254;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2452__delay_2451__delay_2450___cond_2177 <= __delay_data_2451__delay_2450__delay_2449___cond_2177;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2469__delay_2468__delay_2467___cond_2184 <= __delay_data_2468__delay_2467__delay_2466___cond_2184;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2486__delay_2485__delay_2484___plus_2245 <= __delay_data_2485__delay_2484__delay_2483___plus_2245;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2504__delay_2503__delay_2502__delay_2501___eq_2251 <= __delay_data_2503__delay_2502__delay_2501__delay_2500___eq_2251;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2533__delay_2532__delay_2531__delay_2530___eq_2254 <= __delay_data_2532__delay_2531__delay_2530__delay_2529___eq_2254;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2453__delay_2452__delay_2451___cond_2177 <= __delay_data_2452__delay_2451__delay_2450___cond_2177;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2470__delay_2469__delay_2468___cond_2184 <= __delay_data_2469__delay_2468__delay_2467___cond_2184;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2487__delay_2486__delay_2485___plus_2245 <= __delay_data_2486__delay_2485__delay_2484___plus_2245;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2505__delay_2504__delay_2503__delay_2502___eq_2251 <= __delay_data_2504__delay_2503__delay_2502__delay_2501___eq_2251;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2534__delay_2533__delay_2532__delay_2531___eq_2254 <= __delay_data_2533__delay_2532__delay_2531__delay_2530___eq_2254;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2454__delay_2453__delay_2452___cond_2177 <= __delay_data_2453__delay_2452__delay_2451___cond_2177;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2471__delay_2470__delay_2469___cond_2184 <= __delay_data_2470__delay_2469__delay_2468___cond_2184;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2488__delay_2487__delay_2486___plus_2245 <= __delay_data_2487__delay_2486__delay_2485___plus_2245;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2506__delay_2505__delay_2504__delay_2503___eq_2251 <= __delay_data_2505__delay_2504__delay_2503__delay_2502___eq_2251;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2535__delay_2534__delay_2533__delay_2532___eq_2254 <= __delay_data_2534__delay_2533__delay_2532__delay_2531___eq_2254;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _plus_data_2243 <= __substreamoutput_data_2241 + __delay_data_2454__delay_2453__delay_2452___cond_2177;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2472__delay_2471__delay_2470___cond_2184 <= __delay_data_2471__delay_2470__delay_2469___cond_2184;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2489__delay_2488__delay_2487___plus_2245 <= __delay_data_2488__delay_2487__delay_2486___plus_2245;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2507__delay_2506__delay_2505__delay_2504___eq_2251 <= __delay_data_2506__delay_2505__delay_2504__delay_2503___eq_2251;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2536__delay_2535__delay_2534__delay_2533___eq_2254 <= __delay_data_2535__delay_2534__delay_2533__delay_2532___eq_2254;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2548__substreamoutput_2242 <= __substreamoutput_data_2242;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2508__delay_2507__delay_2506__delay_2505___eq_2251 <= __delay_data_2507__delay_2506__delay_2505__delay_2504___eq_2251;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2537__delay_2536__delay_2535__delay_2534___eq_2254 <= __delay_data_2536__delay_2535__delay_2534__delay_2533___eq_2254;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2549__delay_2548__substreamoutput_2242 <= __delay_data_2548__substreamoutput_2242;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2509__delay_2508__delay_2507__delay_2506___eq_2251 <= __delay_data_2508__delay_2507__delay_2506__delay_2505___eq_2251;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2538__delay_2537__delay_2536__delay_2535___eq_2254 <= __delay_data_2537__delay_2536__delay_2535__delay_2534___eq_2254;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2550__delay_2549____substreamoutput_2242 <= __delay_data_2549__delay_2548__substreamoutput_2242;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2510__delay_2509__delay_2508__delay_2507___eq_2251 <= __delay_data_2509__delay_2508__delay_2507__delay_2506___eq_2251;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2539__delay_2538__delay_2537__delay_2536___eq_2254 <= __delay_data_2538__delay_2537__delay_2536__delay_2535___eq_2254;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2551__delay_2550____substreamoutput_2242 <= __delay_data_2550__delay_2549____substreamoutput_2242;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2511__delay_2510__delay_2509__delay_2508___eq_2251 <= __delay_data_2510__delay_2509__delay_2508__delay_2507___eq_2251;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2540__delay_2539__delay_2538__delay_2537___eq_2254 <= __delay_data_2539__delay_2538__delay_2537__delay_2536___eq_2254;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2552__delay_2551____substreamoutput_2242 <= __delay_data_2551__delay_2550____substreamoutput_2242;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2512__delay_2511__delay_2510__delay_2509___eq_2251 <= __delay_data_2511__delay_2510__delay_2509__delay_2508___eq_2251;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2541__delay_2540__delay_2539__delay_2538___eq_2254 <= __delay_data_2540__delay_2539__delay_2538__delay_2537___eq_2254;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2553__delay_2552____substreamoutput_2242 <= __delay_data_2552__delay_2551____substreamoutput_2242;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2513__delay_2512__delay_2511__delay_2510___eq_2251 <= __delay_data_2512__delay_2511__delay_2510__delay_2509___eq_2251;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2542__delay_2541__delay_2540__delay_2539___eq_2254 <= __delay_data_2541__delay_2540__delay_2539__delay_2538___eq_2254;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2554__delay_2553____substreamoutput_2242 <= __delay_data_2553__delay_2552____substreamoutput_2242;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2514__delay_2513__delay_2512__delay_2511___eq_2251 <= __delay_data_2513__delay_2512__delay_2511__delay_2510___eq_2251;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2543__delay_2542__delay_2541__delay_2540___eq_2254 <= __delay_data_2542__delay_2541__delay_2540__delay_2539___eq_2254;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2555__delay_2554____substreamoutput_2242 <= __delay_data_2554__delay_2553____substreamoutput_2242;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2515__delay_2514__delay_2513__delay_2512___eq_2251 <= __delay_data_2514__delay_2513__delay_2512__delay_2511___eq_2251;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2544__delay_2543__delay_2542__delay_2541___eq_2254 <= __delay_data_2543__delay_2542__delay_2541__delay_2540___eq_2254;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2556__delay_2555____substreamoutput_2242 <= __delay_data_2555__delay_2554____substreamoutput_2242;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2516__delay_2515__delay_2514__delay_2513___eq_2251 <= __delay_data_2515__delay_2514__delay_2513__delay_2512___eq_2251;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2545__delay_2544__delay_2543__delay_2542___eq_2254 <= __delay_data_2544__delay_2543__delay_2542__delay_2541___eq_2254;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2557__delay_2556____substreamoutput_2242 <= __delay_data_2556__delay_2555____substreamoutput_2242;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _greaterthan_data_2248 <= __substreamoutput_data_2246 > 1'sd0;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2490__substreamoutput_2246 <= __substreamoutput_data_2246;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2517__delay_2516__delay_2515__delay_2514___eq_2251 <= __delay_data_2516__delay_2515__delay_2514__delay_2513___eq_2251;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2546__delay_2545__delay_2544__delay_2543___eq_2254 <= __delay_data_2545__delay_2544__delay_2543__delay_2542___eq_2254;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2558__delay_2557____substreamoutput_2242 <= __delay_data_2557__delay_2556____substreamoutput_2242;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _cond_data_2250 <= (_greaterthan_data_2248)? __delay_data_2490__substreamoutput_2246 : 1'sd0;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2518__delay_2517__delay_2516__delay_2515___eq_2251 <= __delay_data_2517__delay_2516__delay_2515__delay_2514___eq_2251;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2519__delay_2490__substreamoutput_2246 <= __delay_data_2490__substreamoutput_2246;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2547__delay_2546__delay_2545__delay_2544___eq_2254 <= __delay_data_2546__delay_2545__delay_2544__delay_2543___eq_2254;
      end 
      if(_stream_matmul_11_stream_oready) begin
        __delay_data_2559__delay_2558____substreamoutput_2242 <= __delay_data_2558__delay_2557____substreamoutput_2242;
      end 
      if(_set_flag_1356) begin
        _stream_matmul_11_parameter_0_next_parameter_data <= cparam_matmul_11_stream_reduce_size;
      end 
      if(_stream_matmul_11_source_start) begin
        __variable_wdata_2156 <= _stream_matmul_11_parameter_0_next_parameter_data;
      end 
      if(_set_flag_1357) begin
        _stream_matmul_11_parameter_1_next_parameter_data <= matmul_11_col_select;
      end 
      if(_stream_matmul_11_source_start) begin
        __variable_wdata_2157 <= _stream_matmul_11_parameter_1_next_parameter_data;
      end 
      if(_set_flag_1358) begin
        _stream_matmul_11_parameter_2_next_parameter_data <= matmul_11_row_select_buf;
      end 
      if(_stream_matmul_11_source_start) begin
        __variable_wdata_2158 <= _stream_matmul_11_parameter_2_next_parameter_data;
      end 
      if(_set_flag_1359) begin
        _stream_matmul_11_parameter_3_next_parameter_data <= matmul_11_stream_pad_masks;
      end 
      if(_stream_matmul_11_source_start) begin
        __variable_wdata_2159 <= _stream_matmul_11_parameter_3_next_parameter_data;
      end 
      if(_set_flag_1360) begin
        _stream_matmul_11_parameter_4_next_parameter_data <= cparam_matmul_11_stream_omit_mask;
      end 
      if(_stream_matmul_11_source_start) begin
        __variable_wdata_2160 <= _stream_matmul_11_parameter_4_next_parameter_data;
      end 
      if(_set_flag_1361) begin
        _stream_matmul_11_parameter_6_next_parameter_data <= cparam_matmul_11_bias_scala;
      end 
      if(_stream_matmul_11_source_start) begin
        __variable_wdata_2171 <= _stream_matmul_11_parameter_6_next_parameter_data;
      end 
      if(_set_flag_1362) begin
        _stream_matmul_11_source_7_source_mode <= 5'b10;
        _stream_matmul_11_source_7_source_offset <= (cparam_matmul_11_bias_num == 1)? 0 : matmul_11_och_count_buf;
      end 
      if(_set_flag_1362) begin
        _source_stream_matmul_11_source_7_pat_size_0 <= cparam_matmul_11_stream_reduce_size;
        _source_stream_matmul_11_source_7_pat_stride_0 <= 0;
      end 
      if(_set_flag_1362) begin
        _source_stream_matmul_11_source_7_pat_size_1 <= matmul_11_next_stream_num_ops;
        _source_stream_matmul_11_source_7_pat_stride_1 <= (cparam_matmul_11_bias_num == 1)? 0 : 1;
      end 
      if(_set_flag_1362) begin
        _source_stream_matmul_11_source_7_pat_size_2 <= 1;
        _source_stream_matmul_11_source_7_pat_stride_2 <= 0;
      end 
      if(_set_flag_1362) begin
        _source_stream_matmul_11_source_7_pat_size_3 <= 1;
        _source_stream_matmul_11_source_7_pat_stride_3 <= 0;
      end 
      if(_set_flag_1362) begin
        _stream_matmul_11_source_7_source_sel <= 1;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_7_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _stream_matmul_11_source_7_source_offset_buf <= _stream_matmul_11_source_7_source_offset;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_7_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_7_pat_cur_offset_0 <= 0;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_7_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_7_pat_cur_offset_1 <= 0;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_7_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_7_pat_cur_offset_2 <= 0;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_7_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_7_pat_cur_offset_3 <= 0;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_7_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_7_pat_count_0 <= _source_stream_matmul_11_source_7_pat_size_0 - 1;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_7_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_7_pat_count_1 <= _source_stream_matmul_11_source_7_pat_size_1 - 1;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_7_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_7_pat_count_2 <= _source_stream_matmul_11_source_7_pat_size_2 - 1;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_7_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_7_pat_count_3 <= _source_stream_matmul_11_source_7_pat_size_3 - 1;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_7_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_7_pat_size_buf_0 <= _source_stream_matmul_11_source_7_pat_size_0;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_7_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_7_pat_size_buf_1 <= _source_stream_matmul_11_source_7_pat_size_1;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_7_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_7_pat_size_buf_2 <= _source_stream_matmul_11_source_7_pat_size_2;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_7_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_7_pat_size_buf_3 <= _source_stream_matmul_11_source_7_pat_size_3;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_7_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_7_pat_stride_buf_0 <= _source_stream_matmul_11_source_7_pat_stride_0;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_7_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_7_pat_stride_buf_1 <= _source_stream_matmul_11_source_7_pat_stride_1;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_7_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_7_pat_stride_buf_2 <= _source_stream_matmul_11_source_7_pat_stride_2;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_7_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_7_pat_stride_buf_3 <= _source_stream_matmul_11_source_7_pat_stride_3;
      end 
      if(_stream_matmul_11_stream_oready && _stream_matmul_11_source_busy && _stream_matmul_11_is_root) begin
        __variable_wdata_2172 <= _stream_matmul_11_source_7_source_ram_rdata;
      end 
      if((_stream_matmul_11_source_7_source_pat_fsm_0 == 1) && _stream_matmul_11_stream_oready) begin
        _stream_matmul_11_source_7_idle <= 0;
        _stream_matmul_11_source_7_source_ram_raddr <= _stream_matmul_11_source_7_source_pat_all_offset;
        _stream_matmul_11_source_7_source_ram_renable <= 1;
      end 
      if((_stream_matmul_11_source_7_source_pat_fsm_0 == 1) && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_7_pat_cur_offset_0 <= _source_stream_matmul_11_source_7_pat_cur_offset_0 + _source_stream_matmul_11_source_7_pat_stride_buf_0;
        _source_stream_matmul_11_source_7_pat_count_0 <= _source_stream_matmul_11_source_7_pat_count_0 - 1;
      end 
      if((_stream_matmul_11_source_7_source_pat_fsm_0 == 1) && (_source_stream_matmul_11_source_7_pat_count_0 == 0) && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_7_pat_cur_offset_0 <= 0;
        _source_stream_matmul_11_source_7_pat_count_0 <= _source_stream_matmul_11_source_7_pat_size_buf_0 - 1;
      end 
      if((_stream_matmul_11_source_7_source_pat_fsm_0 == 1) && (_source_stream_matmul_11_source_7_pat_count_0 == 0) && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_7_pat_cur_offset_1 <= _source_stream_matmul_11_source_7_pat_cur_offset_1 + _source_stream_matmul_11_source_7_pat_stride_buf_1;
        _source_stream_matmul_11_source_7_pat_count_1 <= _source_stream_matmul_11_source_7_pat_count_1 - 1;
      end 
      if((_stream_matmul_11_source_7_source_pat_fsm_0 == 1) && (_source_stream_matmul_11_source_7_pat_count_0 == 0) && (_source_stream_matmul_11_source_7_pat_count_1 == 0) && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_7_pat_cur_offset_1 <= 0;
        _source_stream_matmul_11_source_7_pat_count_1 <= _source_stream_matmul_11_source_7_pat_size_buf_1 - 1;
      end 
      if((_stream_matmul_11_source_7_source_pat_fsm_0 == 1) && ((_source_stream_matmul_11_source_7_pat_count_0 == 0) && (_source_stream_matmul_11_source_7_pat_count_1 == 0)) && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_7_pat_cur_offset_2 <= _source_stream_matmul_11_source_7_pat_cur_offset_2 + _source_stream_matmul_11_source_7_pat_stride_buf_2;
        _source_stream_matmul_11_source_7_pat_count_2 <= _source_stream_matmul_11_source_7_pat_count_2 - 1;
      end 
      if((_stream_matmul_11_source_7_source_pat_fsm_0 == 1) && ((_source_stream_matmul_11_source_7_pat_count_0 == 0) && (_source_stream_matmul_11_source_7_pat_count_1 == 0)) && (_source_stream_matmul_11_source_7_pat_count_2 == 0) && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_7_pat_cur_offset_2 <= 0;
        _source_stream_matmul_11_source_7_pat_count_2 <= _source_stream_matmul_11_source_7_pat_size_buf_2 - 1;
      end 
      if((_stream_matmul_11_source_7_source_pat_fsm_0 == 1) && ((_source_stream_matmul_11_source_7_pat_count_0 == 0) && (_source_stream_matmul_11_source_7_pat_count_1 == 0) && (_source_stream_matmul_11_source_7_pat_count_2 == 0)) && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_7_pat_cur_offset_3 <= _source_stream_matmul_11_source_7_pat_cur_offset_3 + _source_stream_matmul_11_source_7_pat_stride_buf_3;
        _source_stream_matmul_11_source_7_pat_count_3 <= _source_stream_matmul_11_source_7_pat_count_3 - 1;
      end 
      if((_stream_matmul_11_source_7_source_pat_fsm_0 == 1) && ((_source_stream_matmul_11_source_7_pat_count_0 == 0) && (_source_stream_matmul_11_source_7_pat_count_1 == 0) && (_source_stream_matmul_11_source_7_pat_count_2 == 0)) && (_source_stream_matmul_11_source_7_pat_count_3 == 0) && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_7_pat_cur_offset_3 <= 0;
        _source_stream_matmul_11_source_7_pat_count_3 <= _source_stream_matmul_11_source_7_pat_size_buf_3 - 1;
      end 
      if((_stream_matmul_11_source_7_source_pat_fsm_0 == 1) && _stream_matmul_11_source_stop && _stream_matmul_11_stream_oready) begin
        _stream_matmul_11_source_7_source_ram_renable <= 0;
        _stream_matmul_11_source_7_idle <= 1;
      end 
      if((_stream_matmul_11_source_7_source_pat_fsm_0 == 2) && _stream_matmul_11_stream_oready) begin
        _stream_matmul_11_source_7_source_ram_renable <= 0;
        _stream_matmul_11_source_7_idle <= 1;
      end 
      if(_set_flag_1371) begin
        _stream_matmul_11_parameter_8_next_parameter_data <= cparam_matmul_11_scale_scala;
      end 
      if(_stream_matmul_11_source_start) begin
        __variable_wdata_2178 <= _stream_matmul_11_parameter_8_next_parameter_data;
      end 
      if(_set_flag_1372) begin
        _stream_matmul_11_source_9_source_mode <= 5'b10;
        _stream_matmul_11_source_9_source_offset <= (cparam_matmul_11_scale_num == 1)? 0 : matmul_11_och_count_buf;
      end 
      if(_set_flag_1372) begin
        _source_stream_matmul_11_source_9_pat_size_0 <= cparam_matmul_11_stream_reduce_size;
        _source_stream_matmul_11_source_9_pat_stride_0 <= 0;
      end 
      if(_set_flag_1372) begin
        _source_stream_matmul_11_source_9_pat_size_1 <= matmul_11_next_stream_num_ops;
        _source_stream_matmul_11_source_9_pat_stride_1 <= (cparam_matmul_11_scale_num == 1)? 0 : 1;
      end 
      if(_set_flag_1372) begin
        _source_stream_matmul_11_source_9_pat_size_2 <= 1;
        _source_stream_matmul_11_source_9_pat_stride_2 <= 0;
      end 
      if(_set_flag_1372) begin
        _source_stream_matmul_11_source_9_pat_size_3 <= 1;
        _source_stream_matmul_11_source_9_pat_stride_3 <= 0;
      end 
      if(_set_flag_1372) begin
        _stream_matmul_11_source_9_source_sel <= 2;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_9_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _stream_matmul_11_source_9_source_offset_buf <= _stream_matmul_11_source_9_source_offset;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_9_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_9_pat_cur_offset_0 <= 0;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_9_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_9_pat_cur_offset_1 <= 0;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_9_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_9_pat_cur_offset_2 <= 0;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_9_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_9_pat_cur_offset_3 <= 0;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_9_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_9_pat_count_0 <= _source_stream_matmul_11_source_9_pat_size_0 - 1;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_9_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_9_pat_count_1 <= _source_stream_matmul_11_source_9_pat_size_1 - 1;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_9_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_9_pat_count_2 <= _source_stream_matmul_11_source_9_pat_size_2 - 1;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_9_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_9_pat_count_3 <= _source_stream_matmul_11_source_9_pat_size_3 - 1;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_9_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_9_pat_size_buf_0 <= _source_stream_matmul_11_source_9_pat_size_0;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_9_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_9_pat_size_buf_1 <= _source_stream_matmul_11_source_9_pat_size_1;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_9_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_9_pat_size_buf_2 <= _source_stream_matmul_11_source_9_pat_size_2;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_9_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_9_pat_size_buf_3 <= _source_stream_matmul_11_source_9_pat_size_3;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_9_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_9_pat_stride_buf_0 <= _source_stream_matmul_11_source_9_pat_stride_0;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_9_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_9_pat_stride_buf_1 <= _source_stream_matmul_11_source_9_pat_stride_1;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_9_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_9_pat_stride_buf_2 <= _source_stream_matmul_11_source_9_pat_stride_2;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_9_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_9_pat_stride_buf_3 <= _source_stream_matmul_11_source_9_pat_stride_3;
      end 
      if(_stream_matmul_11_stream_oready && _stream_matmul_11_source_busy && _stream_matmul_11_is_root) begin
        __variable_wdata_2179 <= _stream_matmul_11_source_9_source_ram_rdata;
      end 
      if((_stream_matmul_11_source_9_source_pat_fsm_1 == 1) && _stream_matmul_11_stream_oready) begin
        _stream_matmul_11_source_9_idle <= 0;
        _stream_matmul_11_source_9_source_ram_raddr <= _stream_matmul_11_source_9_source_pat_all_offset;
        _stream_matmul_11_source_9_source_ram_renable <= 1;
      end 
      if((_stream_matmul_11_source_9_source_pat_fsm_1 == 1) && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_9_pat_cur_offset_0 <= _source_stream_matmul_11_source_9_pat_cur_offset_0 + _source_stream_matmul_11_source_9_pat_stride_buf_0;
        _source_stream_matmul_11_source_9_pat_count_0 <= _source_stream_matmul_11_source_9_pat_count_0 - 1;
      end 
      if((_stream_matmul_11_source_9_source_pat_fsm_1 == 1) && (_source_stream_matmul_11_source_9_pat_count_0 == 0) && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_9_pat_cur_offset_0 <= 0;
        _source_stream_matmul_11_source_9_pat_count_0 <= _source_stream_matmul_11_source_9_pat_size_buf_0 - 1;
      end 
      if((_stream_matmul_11_source_9_source_pat_fsm_1 == 1) && (_source_stream_matmul_11_source_9_pat_count_0 == 0) && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_9_pat_cur_offset_1 <= _source_stream_matmul_11_source_9_pat_cur_offset_1 + _source_stream_matmul_11_source_9_pat_stride_buf_1;
        _source_stream_matmul_11_source_9_pat_count_1 <= _source_stream_matmul_11_source_9_pat_count_1 - 1;
      end 
      if((_stream_matmul_11_source_9_source_pat_fsm_1 == 1) && (_source_stream_matmul_11_source_9_pat_count_0 == 0) && (_source_stream_matmul_11_source_9_pat_count_1 == 0) && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_9_pat_cur_offset_1 <= 0;
        _source_stream_matmul_11_source_9_pat_count_1 <= _source_stream_matmul_11_source_9_pat_size_buf_1 - 1;
      end 
      if((_stream_matmul_11_source_9_source_pat_fsm_1 == 1) && ((_source_stream_matmul_11_source_9_pat_count_0 == 0) && (_source_stream_matmul_11_source_9_pat_count_1 == 0)) && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_9_pat_cur_offset_2 <= _source_stream_matmul_11_source_9_pat_cur_offset_2 + _source_stream_matmul_11_source_9_pat_stride_buf_2;
        _source_stream_matmul_11_source_9_pat_count_2 <= _source_stream_matmul_11_source_9_pat_count_2 - 1;
      end 
      if((_stream_matmul_11_source_9_source_pat_fsm_1 == 1) && ((_source_stream_matmul_11_source_9_pat_count_0 == 0) && (_source_stream_matmul_11_source_9_pat_count_1 == 0)) && (_source_stream_matmul_11_source_9_pat_count_2 == 0) && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_9_pat_cur_offset_2 <= 0;
        _source_stream_matmul_11_source_9_pat_count_2 <= _source_stream_matmul_11_source_9_pat_size_buf_2 - 1;
      end 
      if((_stream_matmul_11_source_9_source_pat_fsm_1 == 1) && ((_source_stream_matmul_11_source_9_pat_count_0 == 0) && (_source_stream_matmul_11_source_9_pat_count_1 == 0) && (_source_stream_matmul_11_source_9_pat_count_2 == 0)) && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_9_pat_cur_offset_3 <= _source_stream_matmul_11_source_9_pat_cur_offset_3 + _source_stream_matmul_11_source_9_pat_stride_buf_3;
        _source_stream_matmul_11_source_9_pat_count_3 <= _source_stream_matmul_11_source_9_pat_count_3 - 1;
      end 
      if((_stream_matmul_11_source_9_source_pat_fsm_1 == 1) && ((_source_stream_matmul_11_source_9_pat_count_0 == 0) && (_source_stream_matmul_11_source_9_pat_count_1 == 0) && (_source_stream_matmul_11_source_9_pat_count_2 == 0)) && (_source_stream_matmul_11_source_9_pat_count_3 == 0) && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_9_pat_cur_offset_3 <= 0;
        _source_stream_matmul_11_source_9_pat_count_3 <= _source_stream_matmul_11_source_9_pat_size_buf_3 - 1;
      end 
      if((_stream_matmul_11_source_9_source_pat_fsm_1 == 1) && _stream_matmul_11_source_stop && _stream_matmul_11_stream_oready) begin
        _stream_matmul_11_source_9_source_ram_renable <= 0;
        _stream_matmul_11_source_9_idle <= 1;
      end 
      if((_stream_matmul_11_source_9_source_pat_fsm_1 == 2) && _stream_matmul_11_stream_oready) begin
        _stream_matmul_11_source_9_source_ram_renable <= 0;
        _stream_matmul_11_source_9_idle <= 1;
      end 
      if(_set_flag_1381) begin
        _stream_matmul_11_parameter_10_next_parameter_data <= 1;
      end 
      if(_stream_matmul_11_source_start) begin
        __variable_wdata_2185 <= _stream_matmul_11_parameter_10_next_parameter_data;
      end 
      if(_set_flag_1382) begin
        _stream_matmul_11_source_11_source_mode <= 5'b0;
        _stream_matmul_11_source_11_source_empty_data <= 0;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_stream_oready && !(|(_stream_matmul_11_source_11_source_mode & 5'b0))) begin
        _stream_matmul_11_source_11_idle <= 1;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_stream_oready && !(|(_stream_matmul_11_source_11_source_mode & 5'b0)) && _stream_matmul_11_is_root) begin
        __variable_wdata_2186 <= _stream_matmul_11_source_11_source_empty_data;
      end 
      if(_set_flag_1383) begin
        _stream_matmul_11_parameter_12_next_parameter_data <= 1;
      end 
      if(_stream_matmul_11_source_start) begin
        __variable_wdata_2192 <= _stream_matmul_11_parameter_12_next_parameter_data;
      end 
      if(_set_flag_1384) begin
        _stream_matmul_11_source_13_source_mode <= 5'b0;
        _stream_matmul_11_source_13_source_empty_data <= 0;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_stream_oready && !(|(_stream_matmul_11_source_13_source_mode & 5'b0))) begin
        _stream_matmul_11_source_13_idle <= 1;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_stream_oready && !(|(_stream_matmul_11_source_13_source_mode & 5'b0)) && _stream_matmul_11_is_root) begin
        __variable_wdata_2193 <= _stream_matmul_11_source_13_source_empty_data;
      end 
      if(_set_flag_1385) begin
        _stream_matmul_11_parameter_14_next_parameter_data <= 1;
      end 
      if(_stream_matmul_11_source_start) begin
        __variable_wdata_2199 <= _stream_matmul_11_parameter_14_next_parameter_data;
      end 
      if(_set_flag_1386) begin
        _stream_matmul_11_source_15_source_mode <= 5'b0;
        _stream_matmul_11_source_15_source_empty_data <= 0;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_stream_oready && !(|(_stream_matmul_11_source_15_source_mode & 5'b0))) begin
        _stream_matmul_11_source_15_idle <= 1;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_stream_oready && !(|(_stream_matmul_11_source_15_source_mode & 5'b0)) && _stream_matmul_11_is_root) begin
        __variable_wdata_2200 <= _stream_matmul_11_source_15_source_empty_data;
      end 
      if(_set_flag_1387) begin
        _stream_matmul_11_parameter_16_next_parameter_data <= cparam_matmul_11_cshamt_mul_value;
      end 
      if(_stream_matmul_11_source_start) begin
        __variable_wdata_2206 <= _stream_matmul_11_parameter_16_next_parameter_data;
      end 
      if(_set_flag_1388) begin
        _stream_matmul_11_parameter_17_next_parameter_data <= cparam_matmul_11_cshamt_sum_value;
      end 
      if(_stream_matmul_11_source_start) begin
        __variable_wdata_2207 <= _stream_matmul_11_parameter_17_next_parameter_data;
      end 
      if(_set_flag_1389) begin
        _stream_matmul_11_parameter_18_next_parameter_data <= cparam_matmul_11_cshamt_out_value;
      end 
      if(_stream_matmul_11_source_start) begin
        __variable_wdata_2208 <= _stream_matmul_11_parameter_18_next_parameter_data;
      end 
      if(_set_flag_1390) begin
        _stream_matmul_11_parameter_19_next_parameter_data <= cparam_matmul_11_act_func_index;
      end 
      if(_stream_matmul_11_source_start) begin
        __variable_wdata_2209 <= _stream_matmul_11_parameter_19_next_parameter_data;
      end 
      if(_set_flag_1391) begin
        _stream_matmul_11_source_20_source_mode <= 5'b10;
        _stream_matmul_11_source_20_source_offset <= matmul_11_stream_act_local_0 + matmul_11_act_page_comp_offset_buf_0;
      end 
      if(_set_flag_1391) begin
        _source_stream_matmul_11_source_20_pat_size_0 <= cparam_matmul_11_stream_reduce_size;
        _source_stream_matmul_11_source_20_pat_stride_0 <= 1;
      end 
      if(_set_flag_1391) begin
        _source_stream_matmul_11_source_20_pat_size_1 <= matmul_11_next_stream_num_ops;
        _source_stream_matmul_11_source_20_pat_stride_1 <= 0;
      end 
      if(_set_flag_1391) begin
        _source_stream_matmul_11_source_20_pat_size_2 <= 1;
        _source_stream_matmul_11_source_20_pat_stride_2 <= 0;
      end 
      if(_set_flag_1391) begin
        _source_stream_matmul_11_source_20_pat_size_3 <= 1;
        _source_stream_matmul_11_source_20_pat_stride_3 <= 0;
      end 
      if(_set_flag_1391) begin
        _stream_matmul_11_source_20_source_sel <= 3;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_20_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _stream_matmul_11_source_20_source_offset_buf <= _stream_matmul_11_source_20_source_offset;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_20_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_20_pat_cur_offset_0 <= 0;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_20_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_20_pat_cur_offset_1 <= 0;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_20_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_20_pat_cur_offset_2 <= 0;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_20_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_20_pat_cur_offset_3 <= 0;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_20_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_20_pat_count_0 <= _source_stream_matmul_11_source_20_pat_size_0 - 1;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_20_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_20_pat_count_1 <= _source_stream_matmul_11_source_20_pat_size_1 - 1;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_20_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_20_pat_count_2 <= _source_stream_matmul_11_source_20_pat_size_2 - 1;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_20_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_20_pat_count_3 <= _source_stream_matmul_11_source_20_pat_size_3 - 1;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_20_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_20_pat_size_buf_0 <= _source_stream_matmul_11_source_20_pat_size_0;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_20_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_20_pat_size_buf_1 <= _source_stream_matmul_11_source_20_pat_size_1;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_20_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_20_pat_size_buf_2 <= _source_stream_matmul_11_source_20_pat_size_2;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_20_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_20_pat_size_buf_3 <= _source_stream_matmul_11_source_20_pat_size_3;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_20_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_20_pat_stride_buf_0 <= _source_stream_matmul_11_source_20_pat_stride_0;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_20_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_20_pat_stride_buf_1 <= _source_stream_matmul_11_source_20_pat_stride_1;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_20_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_20_pat_stride_buf_2 <= _source_stream_matmul_11_source_20_pat_stride_2;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_20_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_20_pat_stride_buf_3 <= _source_stream_matmul_11_source_20_pat_stride_3;
      end 
      if(_stream_matmul_11_stream_oready && _stream_matmul_11_source_busy && _stream_matmul_11_is_root) begin
        __variable_wdata_2210 <= _stream_matmul_11_source_20_source_ram_rdata;
      end 
      if((_stream_matmul_11_source_20_source_pat_fsm_2 == 1) && _stream_matmul_11_stream_oready) begin
        _stream_matmul_11_source_20_idle <= 0;
        _stream_matmul_11_source_20_source_ram_raddr <= _stream_matmul_11_source_20_source_pat_all_offset;
        _stream_matmul_11_source_20_source_ram_renable <= 1;
      end 
      if((_stream_matmul_11_source_20_source_pat_fsm_2 == 1) && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_20_pat_cur_offset_0 <= _source_stream_matmul_11_source_20_pat_cur_offset_0 + _source_stream_matmul_11_source_20_pat_stride_buf_0;
        _source_stream_matmul_11_source_20_pat_count_0 <= _source_stream_matmul_11_source_20_pat_count_0 - 1;
      end 
      if((_stream_matmul_11_source_20_source_pat_fsm_2 == 1) && (_source_stream_matmul_11_source_20_pat_count_0 == 0) && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_20_pat_cur_offset_0 <= 0;
        _source_stream_matmul_11_source_20_pat_count_0 <= _source_stream_matmul_11_source_20_pat_size_buf_0 - 1;
      end 
      if((_stream_matmul_11_source_20_source_pat_fsm_2 == 1) && (_source_stream_matmul_11_source_20_pat_count_0 == 0) && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_20_pat_cur_offset_1 <= _source_stream_matmul_11_source_20_pat_cur_offset_1 + _source_stream_matmul_11_source_20_pat_stride_buf_1;
        _source_stream_matmul_11_source_20_pat_count_1 <= _source_stream_matmul_11_source_20_pat_count_1 - 1;
      end 
      if((_stream_matmul_11_source_20_source_pat_fsm_2 == 1) && (_source_stream_matmul_11_source_20_pat_count_0 == 0) && (_source_stream_matmul_11_source_20_pat_count_1 == 0) && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_20_pat_cur_offset_1 <= 0;
        _source_stream_matmul_11_source_20_pat_count_1 <= _source_stream_matmul_11_source_20_pat_size_buf_1 - 1;
      end 
      if((_stream_matmul_11_source_20_source_pat_fsm_2 == 1) && ((_source_stream_matmul_11_source_20_pat_count_0 == 0) && (_source_stream_matmul_11_source_20_pat_count_1 == 0)) && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_20_pat_cur_offset_2 <= _source_stream_matmul_11_source_20_pat_cur_offset_2 + _source_stream_matmul_11_source_20_pat_stride_buf_2;
        _source_stream_matmul_11_source_20_pat_count_2 <= _source_stream_matmul_11_source_20_pat_count_2 - 1;
      end 
      if((_stream_matmul_11_source_20_source_pat_fsm_2 == 1) && ((_source_stream_matmul_11_source_20_pat_count_0 == 0) && (_source_stream_matmul_11_source_20_pat_count_1 == 0)) && (_source_stream_matmul_11_source_20_pat_count_2 == 0) && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_20_pat_cur_offset_2 <= 0;
        _source_stream_matmul_11_source_20_pat_count_2 <= _source_stream_matmul_11_source_20_pat_size_buf_2 - 1;
      end 
      if((_stream_matmul_11_source_20_source_pat_fsm_2 == 1) && ((_source_stream_matmul_11_source_20_pat_count_0 == 0) && (_source_stream_matmul_11_source_20_pat_count_1 == 0) && (_source_stream_matmul_11_source_20_pat_count_2 == 0)) && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_20_pat_cur_offset_3 <= _source_stream_matmul_11_source_20_pat_cur_offset_3 + _source_stream_matmul_11_source_20_pat_stride_buf_3;
        _source_stream_matmul_11_source_20_pat_count_3 <= _source_stream_matmul_11_source_20_pat_count_3 - 1;
      end 
      if((_stream_matmul_11_source_20_source_pat_fsm_2 == 1) && ((_source_stream_matmul_11_source_20_pat_count_0 == 0) && (_source_stream_matmul_11_source_20_pat_count_1 == 0) && (_source_stream_matmul_11_source_20_pat_count_2 == 0)) && (_source_stream_matmul_11_source_20_pat_count_3 == 0) && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_20_pat_cur_offset_3 <= 0;
        _source_stream_matmul_11_source_20_pat_count_3 <= _source_stream_matmul_11_source_20_pat_size_buf_3 - 1;
      end 
      if((_stream_matmul_11_source_20_source_pat_fsm_2 == 1) && _stream_matmul_11_source_stop && _stream_matmul_11_stream_oready) begin
        _stream_matmul_11_source_20_source_ram_renable <= 0;
        _stream_matmul_11_source_20_idle <= 1;
      end 
      if((_stream_matmul_11_source_20_source_pat_fsm_2 == 2) && _stream_matmul_11_stream_oready) begin
        _stream_matmul_11_source_20_source_ram_renable <= 0;
        _stream_matmul_11_source_20_idle <= 1;
      end 
      if(_set_flag_1400) begin
        _stream_matmul_11_source_21_source_mode <= 5'b10;
        _stream_matmul_11_source_21_source_offset <= matmul_11_filter_page_comp_offset_buf;
      end 
      if(_set_flag_1400) begin
        _source_stream_matmul_11_source_21_pat_size_0 <= cparam_matmul_11_stream_reduce_size;
        _source_stream_matmul_11_source_21_pat_stride_0 <= 1;
      end 
      if(_set_flag_1400) begin
        _source_stream_matmul_11_source_21_pat_size_1 <= matmul_11_next_stream_num_ops;
        _source_stream_matmul_11_source_21_pat_stride_1 <= cparam_matmul_11_stream_aligned_reduce_size;
      end 
      if(_set_flag_1400) begin
        _source_stream_matmul_11_source_21_pat_size_2 <= 1;
        _source_stream_matmul_11_source_21_pat_stride_2 <= 0;
      end 
      if(_set_flag_1400) begin
        _source_stream_matmul_11_source_21_pat_size_3 <= 1;
        _source_stream_matmul_11_source_21_pat_stride_3 <= 0;
      end 
      if(_set_flag_1400) begin
        _stream_matmul_11_source_21_source_sel <= 4;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_21_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _stream_matmul_11_source_21_source_offset_buf <= _stream_matmul_11_source_21_source_offset;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_21_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_21_pat_cur_offset_0 <= 0;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_21_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_21_pat_cur_offset_1 <= 0;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_21_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_21_pat_cur_offset_2 <= 0;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_21_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_21_pat_cur_offset_3 <= 0;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_21_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_21_pat_count_0 <= _source_stream_matmul_11_source_21_pat_size_0 - 1;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_21_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_21_pat_count_1 <= _source_stream_matmul_11_source_21_pat_size_1 - 1;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_21_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_21_pat_count_2 <= _source_stream_matmul_11_source_21_pat_size_2 - 1;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_21_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_21_pat_count_3 <= _source_stream_matmul_11_source_21_pat_size_3 - 1;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_21_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_21_pat_size_buf_0 <= _source_stream_matmul_11_source_21_pat_size_0;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_21_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_21_pat_size_buf_1 <= _source_stream_matmul_11_source_21_pat_size_1;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_21_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_21_pat_size_buf_2 <= _source_stream_matmul_11_source_21_pat_size_2;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_21_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_21_pat_size_buf_3 <= _source_stream_matmul_11_source_21_pat_size_3;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_21_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_21_pat_stride_buf_0 <= _source_stream_matmul_11_source_21_pat_stride_0;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_21_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_21_pat_stride_buf_1 <= _source_stream_matmul_11_source_21_pat_stride_1;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_21_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_21_pat_stride_buf_2 <= _source_stream_matmul_11_source_21_pat_stride_2;
      end 
      if(_stream_matmul_11_source_start && _stream_matmul_11_source_21_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_21_pat_stride_buf_3 <= _source_stream_matmul_11_source_21_pat_stride_3;
      end 
      if(_stream_matmul_11_stream_oready && _stream_matmul_11_source_busy && _stream_matmul_11_is_root) begin
        __variable_wdata_2224 <= _stream_matmul_11_source_21_source_ram_rdata;
      end 
      if((_stream_matmul_11_source_21_source_pat_fsm_3 == 1) && _stream_matmul_11_stream_oready) begin
        _stream_matmul_11_source_21_idle <= 0;
        _stream_matmul_11_source_21_source_ram_raddr <= _stream_matmul_11_source_21_source_pat_all_offset;
        _stream_matmul_11_source_21_source_ram_renable <= 1;
      end 
      if((_stream_matmul_11_source_21_source_pat_fsm_3 == 1) && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_21_pat_cur_offset_0 <= _source_stream_matmul_11_source_21_pat_cur_offset_0 + _source_stream_matmul_11_source_21_pat_stride_buf_0;
        _source_stream_matmul_11_source_21_pat_count_0 <= _source_stream_matmul_11_source_21_pat_count_0 - 1;
      end 
      if((_stream_matmul_11_source_21_source_pat_fsm_3 == 1) && (_source_stream_matmul_11_source_21_pat_count_0 == 0) && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_21_pat_cur_offset_0 <= 0;
        _source_stream_matmul_11_source_21_pat_count_0 <= _source_stream_matmul_11_source_21_pat_size_buf_0 - 1;
      end 
      if((_stream_matmul_11_source_21_source_pat_fsm_3 == 1) && (_source_stream_matmul_11_source_21_pat_count_0 == 0) && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_21_pat_cur_offset_1 <= _source_stream_matmul_11_source_21_pat_cur_offset_1 + _source_stream_matmul_11_source_21_pat_stride_buf_1;
        _source_stream_matmul_11_source_21_pat_count_1 <= _source_stream_matmul_11_source_21_pat_count_1 - 1;
      end 
      if((_stream_matmul_11_source_21_source_pat_fsm_3 == 1) && (_source_stream_matmul_11_source_21_pat_count_0 == 0) && (_source_stream_matmul_11_source_21_pat_count_1 == 0) && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_21_pat_cur_offset_1 <= 0;
        _source_stream_matmul_11_source_21_pat_count_1 <= _source_stream_matmul_11_source_21_pat_size_buf_1 - 1;
      end 
      if((_stream_matmul_11_source_21_source_pat_fsm_3 == 1) && ((_source_stream_matmul_11_source_21_pat_count_0 == 0) && (_source_stream_matmul_11_source_21_pat_count_1 == 0)) && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_21_pat_cur_offset_2 <= _source_stream_matmul_11_source_21_pat_cur_offset_2 + _source_stream_matmul_11_source_21_pat_stride_buf_2;
        _source_stream_matmul_11_source_21_pat_count_2 <= _source_stream_matmul_11_source_21_pat_count_2 - 1;
      end 
      if((_stream_matmul_11_source_21_source_pat_fsm_3 == 1) && ((_source_stream_matmul_11_source_21_pat_count_0 == 0) && (_source_stream_matmul_11_source_21_pat_count_1 == 0)) && (_source_stream_matmul_11_source_21_pat_count_2 == 0) && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_21_pat_cur_offset_2 <= 0;
        _source_stream_matmul_11_source_21_pat_count_2 <= _source_stream_matmul_11_source_21_pat_size_buf_2 - 1;
      end 
      if((_stream_matmul_11_source_21_source_pat_fsm_3 == 1) && ((_source_stream_matmul_11_source_21_pat_count_0 == 0) && (_source_stream_matmul_11_source_21_pat_count_1 == 0) && (_source_stream_matmul_11_source_21_pat_count_2 == 0)) && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_21_pat_cur_offset_3 <= _source_stream_matmul_11_source_21_pat_cur_offset_3 + _source_stream_matmul_11_source_21_pat_stride_buf_3;
        _source_stream_matmul_11_source_21_pat_count_3 <= _source_stream_matmul_11_source_21_pat_count_3 - 1;
      end 
      if((_stream_matmul_11_source_21_source_pat_fsm_3 == 1) && ((_source_stream_matmul_11_source_21_pat_count_0 == 0) && (_source_stream_matmul_11_source_21_pat_count_1 == 0) && (_source_stream_matmul_11_source_21_pat_count_2 == 0)) && (_source_stream_matmul_11_source_21_pat_count_3 == 0) && _stream_matmul_11_stream_oready) begin
        _source_stream_matmul_11_source_21_pat_cur_offset_3 <= 0;
        _source_stream_matmul_11_source_21_pat_count_3 <= _source_stream_matmul_11_source_21_pat_size_buf_3 - 1;
      end 
      if((_stream_matmul_11_source_21_source_pat_fsm_3 == 1) && _stream_matmul_11_source_stop && _stream_matmul_11_stream_oready) begin
        _stream_matmul_11_source_21_source_ram_renable <= 0;
        _stream_matmul_11_source_21_idle <= 1;
      end 
      if((_stream_matmul_11_source_21_source_pat_fsm_3 == 2) && _stream_matmul_11_stream_oready) begin
        _stream_matmul_11_source_21_source_ram_renable <= 0;
        _stream_matmul_11_source_21_idle <= 1;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1410 <= _set_flag_1409;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1411 <= _tmp_1410;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1412 <= _tmp_1411;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1413 <= _tmp_1412;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1414 <= _tmp_1413;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1415 <= _tmp_1414;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1416 <= _tmp_1415;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1417 <= _tmp_1416;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1418 <= _tmp_1417;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1419 <= _tmp_1418;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1420 <= _tmp_1419;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1421 <= _tmp_1420;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1422 <= _tmp_1421;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1423 <= _tmp_1422;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1424 <= _tmp_1423;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1425 <= _tmp_1424;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1426 <= _tmp_1425;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1427 <= _tmp_1426;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1428 <= _tmp_1427;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1429 <= _tmp_1428;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1430 <= _tmp_1429;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1431 <= _tmp_1430;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1432 <= _tmp_1431;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1433 <= _tmp_1432;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1434 <= _tmp_1433;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1435 <= _tmp_1434;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1436 <= _tmp_1435;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1437 <= _tmp_1436;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1438 <= _tmp_1437;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1439 <= _tmp_1438;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1440 <= _tmp_1439;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1443 <= _tmp_1442;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1444 <= _tmp_1443;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1445 <= _tmp_1444;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1446 <= _tmp_1445;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1447 <= _tmp_1446;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1448 <= _tmp_1447;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1449 <= _tmp_1448;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1450 <= _tmp_1449;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1451 <= _tmp_1450;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1452 <= _tmp_1451;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1453 <= _tmp_1452;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1454 <= _tmp_1453;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1455 <= _tmp_1454;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1456 <= _tmp_1455;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1457 <= _tmp_1456;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1458 <= _tmp_1457;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1459 <= _tmp_1458;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1460 <= _tmp_1459;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1461 <= _tmp_1460;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1462 <= _tmp_1461;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1463 <= _tmp_1462;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1464 <= _tmp_1463;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1465 <= _tmp_1464;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1466 <= _tmp_1465;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1467 <= _tmp_1466;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1468 <= _tmp_1467;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1469 <= _tmp_1468;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1470 <= _tmp_1469;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1471 <= _tmp_1470;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1472 <= _tmp_1471;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1473 <= _tmp_1472;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1474 <= matmul_11_next_stream_num_ops;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1475 <= _tmp_1474;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1476 <= _tmp_1475;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1477 <= _tmp_1476;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1478 <= _tmp_1477;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1479 <= _tmp_1478;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1480 <= _tmp_1479;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1481 <= _tmp_1480;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1482 <= _tmp_1481;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1483 <= _tmp_1482;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1484 <= _tmp_1483;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1485 <= _tmp_1484;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1486 <= _tmp_1485;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1487 <= _tmp_1486;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1488 <= _tmp_1487;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1489 <= _tmp_1488;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1490 <= _tmp_1489;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1491 <= _tmp_1490;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1492 <= _tmp_1491;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1493 <= _tmp_1492;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1494 <= _tmp_1493;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1495 <= _tmp_1494;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1496 <= _tmp_1495;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1497 <= _tmp_1496;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1498 <= _tmp_1497;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1499 <= _tmp_1498;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1500 <= _tmp_1499;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1501 <= _tmp_1500;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1502 <= _tmp_1501;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1503 <= _tmp_1502;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1504 <= _tmp_1503;
      end 
      if(_tmp_1440) begin
        _stream_matmul_11_sink_26_sink_mode <= 5'b1;
        _stream_matmul_11_sink_26_sink_offset <= _tmp_1473;
        _stream_matmul_11_sink_26_sink_size <= _tmp_1504;
        _stream_matmul_11_sink_26_sink_stride <= 1;
      end 
      if(_tmp_1440) begin
        _stream_matmul_11_sink_26_sink_sel <= 5;
      end 
      if(_stream_matmul_11_sink_start && _stream_matmul_11_sink_26_sink_mode & 5'b1 && _stream_matmul_11_stream_oready) begin
        _stream_matmul_11_sink_26_sink_offset_buf <= _stream_matmul_11_sink_26_sink_offset;
        _stream_matmul_11_sink_26_sink_size_buf <= _stream_matmul_11_sink_26_sink_size;
        _stream_matmul_11_sink_26_sink_stride_buf <= _stream_matmul_11_sink_26_sink_stride;
      end 
      if((_stream_matmul_11_sink_26_sink_fsm_4 == 1) && _stream_matmul_11_stream_oready) begin
        _stream_matmul_11_sink_26_sink_waddr <= _stream_matmul_11_sink_26_sink_offset_buf - _stream_matmul_11_sink_26_sink_stride_buf;
        _stream_matmul_11_sink_26_sink_count <= _stream_matmul_11_sink_26_sink_size_buf;
      end 
      if((_stream_matmul_11_sink_26_sink_fsm_4 == 2) && stream_matmul_11_sink_27_data && _stream_matmul_11_stream_oready) begin
        _stream_matmul_11_sink_26_sink_waddr <= _stream_matmul_11_sink_26_sink_waddr + _stream_matmul_11_sink_26_sink_stride_buf;
        _stream_matmul_11_sink_26_sink_wdata <= stream_matmul_11_sink_26_data;
        _stream_matmul_11_sink_26_sink_wenable <= 1;
        _stream_matmul_11_sink_26_sink_count <= _stream_matmul_11_sink_26_sink_count - 1;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1517 <= _stream_matmul_11_source_start;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1518 <= _tmp_1517;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1519 <= _tmp_1518;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1520 <= _stream_matmul_11_source_start;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1521 <= _tmp_1520;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1522 <= _tmp_1521;
      end 
      if(_stream_matmul_11_stream_oready && _tmp_1522) begin
        __variable_wdata_2161 <= 1;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1523 <= _stream_matmul_11_source_start;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1524 <= _tmp_1523;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1525 <= _tmp_1524;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1526 <= _tmp_1525;
      end 
      if(_stream_matmul_11_stream_oready && _tmp_1526) begin
        __variable_wdata_2161 <= 0;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1529 <= _tmp_1528;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1532 <= _tmp_1531;
      end 
      if(_stream_matmul_11_stream_oready && _tmp_1532) begin
        __variable_wdata_2161 <= 1;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1533 <= _stream_matmul_11_source_start;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1534 <= _tmp_1533;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1535 <= _tmp_1534;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1536 <= _tmp_1535;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1537 <= _tmp_1536;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1538 <= _tmp_1537;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1539 <= _tmp_1538;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1540 <= _tmp_1539;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1541 <= _tmp_1540;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1542 <= _tmp_1541;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1543 <= _tmp_1542;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1544 <= _tmp_1543;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1545 <= _tmp_1544;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1546 <= _tmp_1545;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1547 <= _tmp_1546;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1548 <= _tmp_1547;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1549 <= _tmp_1548;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1550 <= _tmp_1549;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1551 <= _tmp_1550;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1552 <= _tmp_1551;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1553 <= _tmp_1552;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1554 <= _tmp_1553;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1555 <= _tmp_1554;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1556 <= _tmp_1555;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1557 <= _tmp_1556;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1558 <= _tmp_1557;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1559 <= _tmp_1558;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1560 <= _tmp_1559;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1561 <= _tmp_1560;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1562 <= _tmp_1561;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1563 <= _tmp_1562;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1564 <= _stream_matmul_11_source_stop;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1565 <= _tmp_1564;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1566 <= _tmp_1565;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1567 <= _tmp_1566;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1568 <= _tmp_1567;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1569 <= _tmp_1568;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1570 <= _tmp_1569;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1571 <= _tmp_1570;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1572 <= _tmp_1571;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1573 <= _tmp_1572;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1574 <= _tmp_1573;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1575 <= _tmp_1574;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1576 <= _tmp_1575;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1577 <= _tmp_1576;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1578 <= _tmp_1577;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1579 <= _tmp_1578;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1580 <= _tmp_1579;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1581 <= _tmp_1580;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1582 <= _tmp_1581;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1583 <= _tmp_1582;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1584 <= _tmp_1583;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1585 <= _tmp_1584;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1586 <= _tmp_1585;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1587 <= _tmp_1586;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1588 <= _tmp_1587;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1589 <= _tmp_1588;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1590 <= _tmp_1589;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1591 <= _tmp_1590;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1592 <= _tmp_1591;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1593 <= _tmp_1592;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1594 <= _tmp_1593;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1595 <= _stream_matmul_11_source_busy;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1596 <= _tmp_1595;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1597 <= _tmp_1596;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1598 <= _tmp_1597;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1599 <= _tmp_1598;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1600 <= _tmp_1599;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1601 <= _tmp_1600;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1602 <= _tmp_1601;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1603 <= _tmp_1602;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1604 <= _tmp_1603;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1605 <= _tmp_1604;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1606 <= _tmp_1605;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1607 <= _tmp_1606;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1608 <= _tmp_1607;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1609 <= _tmp_1608;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1610 <= _tmp_1609;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1611 <= _tmp_1610;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1612 <= _tmp_1611;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1613 <= _tmp_1612;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1614 <= _tmp_1613;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1615 <= _tmp_1614;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1616 <= _tmp_1615;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1617 <= _tmp_1616;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1618 <= _tmp_1617;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1619 <= _tmp_1618;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1620 <= _tmp_1619;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1621 <= _tmp_1620;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1622 <= _tmp_1621;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1623 <= _tmp_1622;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1624 <= _tmp_1623;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1625 <= _tmp_1624;
      end 
      if(_stream_matmul_11_stream_oready) begin
        _tmp_1626 <= _stream_matmul_11_sink_busy;
      end 
      if(!_stream_matmul_11_sink_busy && _tmp_1626) begin
        _stream_matmul_11_busy_reg <= 0;
      end 
      if(_stream_matmul_11_source_busy) begin
        _stream_matmul_11_busy_reg <= 1;
      end 
    end
  end

  localparam _stream_matmul_11_fsm_1 = 1;
  localparam _stream_matmul_11_fsm_2 = 2;
  localparam _stream_matmul_11_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_matmul_11_fsm <= _stream_matmul_11_fsm_init;
      _stream_matmul_11_source_start <= 0;
      _stream_matmul_11_source_busy <= 0;
      _stream_matmul_11_stream_ivalid <= 0;
    end else begin
      if(_stream_matmul_11_stream_oready && _tmp_1519) begin
        _stream_matmul_11_stream_ivalid <= 1;
      end 
      if(_stream_matmul_11_stream_oready && _tmp_1529) begin
        _stream_matmul_11_stream_ivalid <= 0;
      end 
      case(_stream_matmul_11_fsm)
        _stream_matmul_11_fsm_init: begin
          if(_stream_matmul_11_run_flag) begin
            _stream_matmul_11_source_start <= 1;
          end 
          if(_stream_matmul_11_run_flag) begin
            _stream_matmul_11_fsm <= _stream_matmul_11_fsm_1;
          end 
        end
        _stream_matmul_11_fsm_1: begin
          if(_stream_matmul_11_source_start && _stream_matmul_11_stream_oready) begin
            _stream_matmul_11_source_start <= 0;
            _stream_matmul_11_source_busy <= 1;
          end 
          if(_stream_matmul_11_source_start && _stream_matmul_11_stream_oready) begin
            _stream_matmul_11_fsm <= _stream_matmul_11_fsm_2;
          end 
        end
        _stream_matmul_11_fsm_2: begin
          if(_stream_matmul_11_stream_oready) begin
            _stream_matmul_11_fsm <= _stream_matmul_11_fsm_3;
          end 
        end
        _stream_matmul_11_fsm_3: begin
          if(_stream_matmul_11_stream_oready && (_stream_matmul_11_source_11_idle && _stream_matmul_11_source_13_idle && _stream_matmul_11_source_15_idle && _stream_matmul_11_source_20_idle && _stream_matmul_11_source_21_idle && _stream_matmul_11_source_7_idle && _stream_matmul_11_source_9_idle && (_stream_matmul_11_fsm == 3))) begin
            _stream_matmul_11_source_busy <= 0;
          end 
          if(_stream_matmul_11_stream_oready && (_stream_matmul_11_source_11_idle && _stream_matmul_11_source_13_idle && _stream_matmul_11_source_15_idle && _stream_matmul_11_source_20_idle && _stream_matmul_11_source_21_idle && _stream_matmul_11_source_7_idle && _stream_matmul_11_source_9_idle && (_stream_matmul_11_fsm == 3)) && _stream_matmul_11_run_flag) begin
            _stream_matmul_11_source_start <= 1;
          end 
          if(_stream_matmul_11_stream_oready && (_stream_matmul_11_source_11_idle && _stream_matmul_11_source_13_idle && _stream_matmul_11_source_15_idle && _stream_matmul_11_source_20_idle && _stream_matmul_11_source_21_idle && _stream_matmul_11_source_7_idle && _stream_matmul_11_source_9_idle && (_stream_matmul_11_fsm == 3))) begin
            _stream_matmul_11_fsm <= _stream_matmul_11_fsm_init;
          end 
          if(_stream_matmul_11_stream_oready && (_stream_matmul_11_source_11_idle && _stream_matmul_11_source_13_idle && _stream_matmul_11_source_15_idle && _stream_matmul_11_source_20_idle && _stream_matmul_11_source_21_idle && _stream_matmul_11_source_7_idle && _stream_matmul_11_source_9_idle && (_stream_matmul_11_fsm == 3)) && _stream_matmul_11_run_flag) begin
            _stream_matmul_11_fsm <= _stream_matmul_11_fsm_1;
          end 
        end
      endcase
    end
  end

  localparam main_fsm_1 = 1;
  localparam main_fsm_2 = 2;
  localparam main_fsm_3 = 3;
  localparam main_fsm_4 = 4;
  localparam main_fsm_5 = 5;
  localparam main_fsm_6 = 6;
  localparam main_fsm_7 = 7;
  localparam main_fsm_8 = 8;
  localparam main_fsm_9 = 9;
  localparam main_fsm_10 = 10;
  localparam main_fsm_11 = 11;
  localparam main_fsm_12 = 12;
  localparam main_fsm_13 = 13;
  localparam main_fsm_14 = 14;
  localparam main_fsm_15 = 15;
  localparam main_fsm_16 = 16;
  localparam main_fsm_17 = 17;
  localparam main_fsm_18 = 18;
  localparam main_fsm_19 = 19;
  localparam main_fsm_20 = 20;
  localparam main_fsm_21 = 21;
  localparam main_fsm_22 = 22;
  localparam main_fsm_23 = 23;
  localparam main_fsm_24 = 24;
  localparam main_fsm_25 = 25;
  localparam main_fsm_26 = 26;
  localparam main_fsm_27 = 27;
  localparam main_fsm_28 = 28;
  localparam main_fsm_29 = 29;
  localparam main_fsm_30 = 30;
  localparam main_fsm_31 = 31;
  localparam main_fsm_32 = 32;
  localparam main_fsm_33 = 33;
  localparam main_fsm_34 = 34;
  localparam main_fsm_35 = 35;
  localparam main_fsm_36 = 36;
  localparam main_fsm_37 = 37;
  localparam main_fsm_38 = 38;
  localparam main_fsm_39 = 39;
  localparam main_fsm_40 = 40;
  localparam main_fsm_41 = 41;
  localparam main_fsm_42 = 42;
  localparam main_fsm_43 = 43;
  localparam main_fsm_44 = 44;
  localparam main_fsm_45 = 45;
  localparam main_fsm_46 = 46;

  always @(posedge CLK) begin
    if(RST) begin
      main_fsm <= main_fsm_init;
      conv2d_4_objaddr <= 0;
      conv2d_4_arg_objaddr_0 <= 0;
      conv2d_4_arg_objaddr_1 <= 0;
      conv2d_4_arg_objaddr_2 <= 0;
      conv2d_4_arg_objaddr_3 <= 0;
      max_pool_serial_6_objaddr <= 0;
      max_pool_serial_6_arg_objaddr_0 <= 0;
      matmul_11_objaddr <= 0;
      matmul_11_arg_objaddr_0 <= 0;
      matmul_11_arg_objaddr_1 <= 0;
      matmul_11_arg_objaddr_2 <= 0;
      matmul_11_arg_objaddr_3 <= 0;
      matmul_11_control_param_index <= 0;
    end else begin
      case(main_fsm)
        main_fsm_init: begin
          if(_saxi_register_4 != 0) begin
            main_fsm <= main_fsm_1;
          end 
        end
        main_fsm_1: begin
          main_fsm <= main_fsm_2;
        end
        main_fsm_2: begin
          main_fsm <= main_fsm_3;
        end
        main_fsm_3: begin
          main_fsm <= main_fsm_4;
        end
        main_fsm_4: begin
          main_fsm <= main_fsm_5;
        end
        main_fsm_5: begin
          conv2d_4_objaddr <= _saxi_register_33;
          main_fsm <= main_fsm_6;
        end
        main_fsm_6: begin
          conv2d_4_arg_objaddr_0 <= _saxi_register_35;
          main_fsm <= main_fsm_7;
        end
        main_fsm_7: begin
          conv2d_4_arg_objaddr_1 <= _saxi_register_36;
          main_fsm <= main_fsm_8;
        end
        main_fsm_8: begin
          conv2d_4_arg_objaddr_2 <= _saxi_register_36 + 1152;
          main_fsm <= main_fsm_9;
        end
        main_fsm_9: begin
          conv2d_4_arg_objaddr_3 <= _saxi_register_36 + 1216;
          main_fsm <= main_fsm_10;
        end
        main_fsm_10: begin
          main_fsm <= main_fsm_11;
        end
        main_fsm_11: begin
          main_fsm <= main_fsm_12;
        end
        main_fsm_12: begin
          if(control_conv2d_4 == 34) begin
            main_fsm <= main_fsm_13;
          end 
        end
        main_fsm_13: begin
          main_fsm <= main_fsm_14;
        end
        main_fsm_14: begin
          max_pool_serial_6_objaddr <= _saxi_register_33 + 50176;
          main_fsm <= main_fsm_15;
        end
        main_fsm_15: begin
          max_pool_serial_6_arg_objaddr_0 <= _saxi_register_33;
          main_fsm <= main_fsm_16;
        end
        main_fsm_16: begin
          main_fsm <= main_fsm_17;
        end
        main_fsm_17: begin
          main_fsm <= main_fsm_18;
        end
        main_fsm_18: begin
          if(control_max_pool_serial_6 == 19) begin
            main_fsm <= main_fsm_19;
          end 
        end
        main_fsm_19: begin
          main_fsm <= main_fsm_20;
        end
        main_fsm_20: begin
          main_fsm <= main_fsm_21;
        end
        main_fsm_21: begin
          main_fsm <= main_fsm_22;
        end
        main_fsm_22: begin
          matmul_11_objaddr <= _saxi_register_33 + 62720;
          main_fsm <= main_fsm_23;
        end
        main_fsm_23: begin
          matmul_11_arg_objaddr_0 <= _saxi_register_33 + 50176;
          main_fsm <= main_fsm_24;
        end
        main_fsm_24: begin
          matmul_11_arg_objaddr_1 <= _saxi_register_36 + 1280;
          main_fsm <= main_fsm_25;
        end
        main_fsm_25: begin
          matmul_11_arg_objaddr_2 <= _saxi_register_36 + 1606912;
          main_fsm <= main_fsm_26;
        end
        main_fsm_26: begin
          matmul_11_arg_objaddr_3 <= _saxi_register_36 + 1607168;
          main_fsm <= main_fsm_27;
        end
        main_fsm_27: begin
          matmul_11_control_param_index <= 0;
          main_fsm <= main_fsm_28;
        end
        main_fsm_28: begin
          main_fsm <= main_fsm_29;
        end
        main_fsm_29: begin
          main_fsm <= main_fsm_30;
        end
        main_fsm_30: begin
          if(control_matmul_11 == 28) begin
            main_fsm <= main_fsm_31;
          end 
        end
        main_fsm_31: begin
          main_fsm <= main_fsm_32;
        end
        main_fsm_32: begin
          matmul_11_objaddr <= _saxi_register_34;
          main_fsm <= main_fsm_33;
        end
        main_fsm_33: begin
          matmul_11_arg_objaddr_0 <= _saxi_register_33 + 62720;
          main_fsm <= main_fsm_34;
        end
        main_fsm_34: begin
          matmul_11_arg_objaddr_1 <= _saxi_register_36 + 1607424;
          main_fsm <= main_fsm_35;
        end
        main_fsm_35: begin
          matmul_11_arg_objaddr_2 <= _saxi_register_36 + 1609984;
          main_fsm <= main_fsm_36;
        end
        main_fsm_36: begin
          matmul_11_arg_objaddr_3 <= _saxi_register_36 + 1610048;
          main_fsm <= main_fsm_37;
        end
        main_fsm_37: begin
          matmul_11_control_param_index <= 1;
          main_fsm <= main_fsm_38;
        end
        main_fsm_38: begin
          main_fsm <= main_fsm_39;
        end
        main_fsm_39: begin
          main_fsm <= main_fsm_40;
        end
        main_fsm_40: begin
          if(control_matmul_11 == 28) begin
            main_fsm <= main_fsm_41;
          end 
        end
        main_fsm_41: begin
          main_fsm <= main_fsm_42;
        end
        main_fsm_42: begin
          main_fsm <= main_fsm_43;
        end
        main_fsm_43: begin
          main_fsm <= main_fsm_44;
        end
        main_fsm_44: begin
          main_fsm <= main_fsm_45;
        end
        main_fsm_45: begin
          main_fsm <= main_fsm_46;
        end
        main_fsm_46: begin
          main_fsm <= main_fsm_init;
        end
      endcase
    end
  end

  localparam control_conv2d_4_1 = 1;
  localparam control_conv2d_4_2 = 2;
  localparam control_conv2d_4_3 = 3;
  localparam control_conv2d_4_4 = 4;
  localparam control_conv2d_4_5 = 5;
  localparam control_conv2d_4_6 = 6;
  localparam control_conv2d_4_7 = 7;
  localparam control_conv2d_4_8 = 8;
  localparam control_conv2d_4_9 = 9;
  localparam control_conv2d_4_10 = 10;
  localparam control_conv2d_4_11 = 11;
  localparam control_conv2d_4_12 = 12;
  localparam control_conv2d_4_13 = 13;
  localparam control_conv2d_4_14 = 14;
  localparam control_conv2d_4_15 = 15;
  localparam control_conv2d_4_16 = 16;
  localparam control_conv2d_4_17 = 17;
  localparam control_conv2d_4_18 = 18;
  localparam control_conv2d_4_19 = 19;
  localparam control_conv2d_4_20 = 20;
  localparam control_conv2d_4_21 = 21;
  localparam control_conv2d_4_22 = 22;
  localparam control_conv2d_4_23 = 23;
  localparam control_conv2d_4_24 = 24;
  localparam control_conv2d_4_25 = 25;
  localparam control_conv2d_4_26 = 26;
  localparam control_conv2d_4_27 = 27;
  localparam control_conv2d_4_28 = 28;
  localparam control_conv2d_4_29 = 29;
  localparam control_conv2d_4_30 = 30;
  localparam control_conv2d_4_31 = 31;
  localparam control_conv2d_4_32 = 32;
  localparam control_conv2d_4_33 = 33;
  localparam control_conv2d_4_34 = 34;

  always @(posedge CLK) begin
    if(RST) begin
      control_conv2d_4 <= control_conv2d_4_init;
      _control_conv2d_4_called <= 0;
      conv2d_4_filter_base_offset <= 0;
      conv2d_4_filter_page_comp_offset <= 0;
      conv2d_4_filter_page_dma_offset <= 0;
      conv2d_4_act_base_offset_row <= 0;
      conv2d_4_act_base_offset_bat <= 0;
      conv2d_4_dma_flag_0 <= 0;
      conv2d_4_dma_flag_1 <= 0;
      conv2d_4_dma_flag_2 <= 0;
      conv2d_4_act_page_comp_offset_0 <= 0;
      conv2d_4_act_page_comp_offset_1 <= 0;
      conv2d_4_act_page_comp_offset_2 <= 0;
      conv2d_4_act_page_dma_offset_0 <= 0;
      conv2d_4_act_page_dma_offset_1 <= 0;
      conv2d_4_act_page_dma_offset_2 <= 0;
      conv2d_4_out_base_offset_val <= 0;
      conv2d_4_out_base_offset_col <= 0;
      conv2d_4_out_base_offset_row <= 0;
      conv2d_4_out_base_offset_bat <= 0;
      conv2d_4_out_base_offset_och <= 0;
      conv2d_4_out_page <= 0;
      conv2d_4_out_page_comp_offset <= 0;
      conv2d_4_out_page_dma_offset <= 0;
      conv2d_4_out_laddr_offset <= 0;
      conv2d_4_sync_out_count <= 0;
      conv2d_4_write_count <= 0;
      conv2d_4_next_out_write_size <= 0;
      conv2d_4_row_count <= 0;
      conv2d_4_bat_count <= 0;
      conv2d_4_och_count <= 0;
      conv2d_4_row_select <= 0;
      conv2d_4_prev_row_count <= 0;
      conv2d_4_prev_bat_count <= 0;
      conv2d_4_prev_och_count <= 0;
      conv2d_4_prev_row_select <= 0;
      conv2d_4_out_col_count <= 0;
      conv2d_4_out_row_count <= 0;
      conv2d_4_out_ram_select <= 0;
      conv2d_4_skip_read_filter <= 0;
      conv2d_4_skip_read_act <= 0;
      conv2d_4_skip_comp <= 0;
      conv2d_4_skip_write_out <= 1;
    end else begin
      case(control_conv2d_4)
        control_conv2d_4_init: begin
          if(main_fsm == 10) begin
            _control_conv2d_4_called <= 1;
          end 
          if(main_fsm == 10) begin
            control_conv2d_4 <= control_conv2d_4_1;
          end 
        end
        control_conv2d_4_1: begin
          control_conv2d_4 <= control_conv2d_4_2;
        end
        control_conv2d_4_2: begin
          conv2d_4_filter_base_offset <= 0;
          conv2d_4_filter_page_comp_offset <= 0;
          conv2d_4_filter_page_dma_offset <= 0;
          conv2d_4_act_base_offset_row <= 0;
          conv2d_4_act_base_offset_bat <= 0;
          conv2d_4_dma_flag_0 <= 1;
          conv2d_4_dma_flag_1 <= 1;
          conv2d_4_dma_flag_2 <= 1;
          conv2d_4_act_page_comp_offset_0 <= 0;
          conv2d_4_act_page_comp_offset_1 <= 0;
          conv2d_4_act_page_comp_offset_2 <= 0;
          conv2d_4_act_page_dma_offset_0 <= 0;
          conv2d_4_act_page_dma_offset_1 <= 0;
          conv2d_4_act_page_dma_offset_2 <= 0;
          conv2d_4_out_base_offset_val <= 0;
          conv2d_4_out_base_offset_col <= 0;
          conv2d_4_out_base_offset_row <= 0;
          conv2d_4_out_base_offset_bat <= 0;
          conv2d_4_out_base_offset_och <= 0;
          conv2d_4_out_page <= 0;
          conv2d_4_out_page_comp_offset <= 0;
          conv2d_4_out_page_dma_offset <= 0;
          conv2d_4_out_laddr_offset <= 0;
          conv2d_4_sync_out_count <= 0;
          conv2d_4_write_count <= 0;
          conv2d_4_next_out_write_size <= (cparam_conv2d_4_max_och_count == 0)? cparam_conv2d_4_out_write_size_res : cparam_conv2d_4_out_write_size;
          conv2d_4_row_count <= 0;
          conv2d_4_bat_count <= 0;
          conv2d_4_och_count <= 0;
          conv2d_4_row_select <= 0;
          conv2d_4_prev_row_count <= 0;
          conv2d_4_prev_bat_count <= 0;
          conv2d_4_prev_och_count <= 0;
          conv2d_4_prev_row_select <= 0;
          conv2d_4_out_col_count <= 0;
          conv2d_4_out_row_count <= 0;
          conv2d_4_out_ram_select <= 0;
          conv2d_4_skip_read_filter <= 0;
          conv2d_4_skip_read_act <= 0;
          conv2d_4_skip_comp <= 0;
          conv2d_4_skip_write_out <= 1;
          if(_maxi_read_req_idle) begin
            control_conv2d_4 <= control_conv2d_4_3;
          end 
        end
        control_conv2d_4_3: begin
          if(_maxi_read_idle) begin
            control_conv2d_4 <= control_conv2d_4_4;
          end 
        end
        control_conv2d_4_4: begin
          if(_maxi_read_req_idle) begin
            control_conv2d_4 <= control_conv2d_4_5;
          end 
        end
        control_conv2d_4_5: begin
          if(_maxi_read_idle) begin
            control_conv2d_4 <= control_conv2d_4_6;
          end 
        end
        control_conv2d_4_6: begin
          if(cparam_conv2d_4_data_stationary == 0) begin
            control_conv2d_4 <= control_conv2d_4_7;
          end 
          if(cparam_conv2d_4_data_stationary == 1) begin
            control_conv2d_4 <= control_conv2d_4_12;
          end 
        end
        control_conv2d_4_7: begin
          control_conv2d_4 <= control_conv2d_4_8;
          if(conv2d_4_skip_read_filter) begin
            control_conv2d_4 <= control_conv2d_4_11;
          end 
        end
        control_conv2d_4_8: begin
          if(_maxi_read_req_idle) begin
            control_conv2d_4 <= control_conv2d_4_9;
          end 
        end
        control_conv2d_4_9: begin
          if(_maxi_read_idle) begin
            control_conv2d_4 <= control_conv2d_4_10;
          end 
        end
        control_conv2d_4_10: begin
          control_conv2d_4 <= control_conv2d_4_11;
        end
        control_conv2d_4_11: begin
          if(cparam_conv2d_4_data_stationary == 0) begin
            control_conv2d_4 <= control_conv2d_4_12;
          end 
          if(cparam_conv2d_4_data_stationary == 1) begin
            control_conv2d_4 <= control_conv2d_4_24;
          end 
        end
        control_conv2d_4_12: begin
          control_conv2d_4 <= control_conv2d_4_13;
          if(conv2d_4_skip_read_act) begin
            control_conv2d_4 <= control_conv2d_4_23;
          end 
        end
        control_conv2d_4_13: begin
          control_conv2d_4 <= control_conv2d_4_14;
          if(conv2d_4_mux_dma_pad_mask_0 || !conv2d_4_mux_dma_flag_0) begin
            control_conv2d_4 <= control_conv2d_4_16;
          end 
        end
        control_conv2d_4_14: begin
          if(_maxi_read_req_idle) begin
            control_conv2d_4 <= control_conv2d_4_15;
          end 
        end
        control_conv2d_4_15: begin
          if(_maxi_read_idle) begin
            control_conv2d_4 <= control_conv2d_4_16;
          end 
        end
        control_conv2d_4_16: begin
          control_conv2d_4 <= control_conv2d_4_17;
          if(conv2d_4_mux_dma_pad_mask_1 || !conv2d_4_mux_dma_flag_1) begin
            control_conv2d_4 <= control_conv2d_4_19;
          end 
        end
        control_conv2d_4_17: begin
          if(_maxi_read_req_idle) begin
            control_conv2d_4 <= control_conv2d_4_18;
          end 
        end
        control_conv2d_4_18: begin
          if(_maxi_read_idle) begin
            control_conv2d_4 <= control_conv2d_4_19;
          end 
        end
        control_conv2d_4_19: begin
          control_conv2d_4 <= control_conv2d_4_20;
          if(conv2d_4_mux_dma_pad_mask_2 || !conv2d_4_mux_dma_flag_2) begin
            control_conv2d_4 <= control_conv2d_4_22;
          end 
        end
        control_conv2d_4_20: begin
          if(_maxi_read_req_idle) begin
            control_conv2d_4 <= control_conv2d_4_21;
          end 
        end
        control_conv2d_4_21: begin
          if(_maxi_read_idle) begin
            control_conv2d_4 <= control_conv2d_4_22;
          end 
        end
        control_conv2d_4_22: begin
          control_conv2d_4 <= control_conv2d_4_23;
        end
        control_conv2d_4_23: begin
          if(cparam_conv2d_4_data_stationary == 0) begin
            control_conv2d_4 <= control_conv2d_4_24;
          end 
          if(cparam_conv2d_4_data_stationary == 1) begin
            control_conv2d_4 <= control_conv2d_4_7;
          end 
        end
        control_conv2d_4_24: begin
          if(_maxi_write_idle) begin
            control_conv2d_4 <= control_conv2d_4_25;
          end 
        end
        control_conv2d_4_25: begin
          if(conv2d_4_comp_fsm == 0) begin
            control_conv2d_4 <= control_conv2d_4_26;
          end 
        end
        control_conv2d_4_26: begin
          control_conv2d_4 <= control_conv2d_4_27;
          if(conv2d_4_skip_write_out) begin
            control_conv2d_4 <= control_conv2d_4_32;
          end 
          if((cparam_conv2d_4_data_stationary == 1) && (conv2d_4_prev_och_count < cparam_conv2d_4_max_och_count)) begin
            control_conv2d_4 <= control_conv2d_4_32;
          end 
        end
        control_conv2d_4_27: begin
          if(conv2d_4_sync_comp_count >= conv2d_4_sync_out_count + cparam_conv2d_4_inc_sync_out) begin
            control_conv2d_4 <= control_conv2d_4_28;
          end 
        end
        control_conv2d_4_28: begin
          if(!conv2d_4_dma_out_mask_0) begin
            control_conv2d_4 <= control_conv2d_4_29;
          end 
          if(conv2d_4_dma_out_mask_0) begin
            control_conv2d_4 <= control_conv2d_4_30;
          end 
        end
        control_conv2d_4_29: begin
          if(_maxi_write_req_idle) begin
            control_conv2d_4 <= control_conv2d_4_30;
          end 
        end
        control_conv2d_4_30: begin
          control_conv2d_4 <= control_conv2d_4_31;
        end
        control_conv2d_4_31: begin
          conv2d_4_write_count <= conv2d_4_write_count + 1;
          if(conv2d_4_out_ram_select == 0) begin
            conv2d_4_out_laddr_offset <= conv2d_4_out_laddr_offset + conv2d_4_next_out_write_size;
          end 
          if((cparam_conv2d_4_data_stationary == 0) && !cparam_conv2d_4_keep_filter) begin
            conv2d_4_out_base_offset_col <= conv2d_4_out_base_offset_col + cparam_conv2d_4_out_col_step;
            conv2d_4_out_col_count <= conv2d_4_out_col_count + 1;
          end 
          conv2d_4_out_ram_select <= conv2d_4_out_ram_select + 1;
          if(conv2d_4_out_ram_select == 0) begin
            conv2d_4_out_ram_select <= 0;
          end 
          conv2d_4_sync_out_count <= conv2d_4_sync_out_count + cparam_conv2d_4_inc_sync_out;
          if((cparam_conv2d_4_data_stationary == 0) && !cparam_conv2d_4_keep_filter && (conv2d_4_write_count >= cparam_conv2d_4_out_num_col - 1) || (cparam_conv2d_4_data_stationary == 0) && cparam_conv2d_4_keep_filter || (cparam_conv2d_4_data_stationary == 1)) begin
            conv2d_4_sync_out_count <= conv2d_4_sync_out_count + (cparam_conv2d_4_inc_sync_out + cparam_conv2d_4_inc_sync_out_res);
          end 
          if((cparam_conv2d_4_data_stationary == 0) && !cparam_conv2d_4_keep_filter) begin
            control_conv2d_4 <= control_conv2d_4_26;
          end 
          if((cparam_conv2d_4_data_stationary == 0) && !cparam_conv2d_4_keep_filter && (conv2d_4_write_count >= cparam_conv2d_4_out_num_col - 1) || (cparam_conv2d_4_data_stationary == 0) && cparam_conv2d_4_keep_filter || (cparam_conv2d_4_data_stationary == 1)) begin
            control_conv2d_4 <= control_conv2d_4_32;
          end 
        end
        control_conv2d_4_32: begin
          if(conv2d_4_update_filter) begin
            conv2d_4_filter_base_offset <= conv2d_4_filter_base_offset + cparam_conv2d_4_filter_base_step;
          end 
          if((cparam_conv2d_4_data_stationary == 1) && (conv2d_4_och_count >= cparam_conv2d_4_max_och_count)) begin
            conv2d_4_filter_base_offset <= 0;
          end 
          if(conv2d_4_update_filter) begin
            conv2d_4_och_count <= conv2d_4_och_count + cparam_conv2d_4_och_count_step;
          end 
          if((cparam_conv2d_4_data_stationary == 1) && (conv2d_4_och_count >= cparam_conv2d_4_max_och_count)) begin
            conv2d_4_och_count <= 0;
          end 
          if(conv2d_4_update_filter) begin
            conv2d_4_filter_page_comp_offset <= conv2d_4_filter_page_comp_offset + cparam_conv2d_4_filter_read_step;
            conv2d_4_filter_page_dma_offset <= conv2d_4_filter_page_dma_offset + cparam_conv2d_4_filter_read_step;
          end 
          if(conv2d_4_update_filter && (conv2d_4_filter_page_comp_offset + cparam_conv2d_4_filter_read_step + cparam_conv2d_4_filter_read_step > 512)) begin
            conv2d_4_filter_page_comp_offset <= 0;
            conv2d_4_filter_page_dma_offset <= 0;
          end 
          if(conv2d_4_update_act) begin
            conv2d_4_act_base_offset_row <= conv2d_4_act_base_offset_row + cparam_conv2d_4_act_row_step;
          end 
          if(conv2d_4_update_act && (conv2d_4_row_count >= cparam_conv2d_4_max_row_count)) begin
            conv2d_4_act_base_offset_row <= 0;
            conv2d_4_act_base_offset_bat <= conv2d_4_act_base_offset_bat + cparam_conv2d_4_act_bat_step;
          end 
          if(conv2d_4_update_act && (conv2d_4_row_count >= cparam_conv2d_4_max_row_count) && (conv2d_4_bat_count >= cparam_conv2d_4_max_bat_count)) begin
            conv2d_4_act_base_offset_bat <= 0;
          end 
          if(!conv2d_4_update_act) begin
            conv2d_4_dma_flag_0 <= 0;
          end 
          if(conv2d_4_update_act) begin
            conv2d_4_dma_flag_0 <= cparam_conv2d_4_dma_flag_conds_0;
          end 
          if(conv2d_4_update_act && (conv2d_4_row_count >= cparam_conv2d_4_max_row_count)) begin
            conv2d_4_dma_flag_0 <= 1;
          end 
          if(!conv2d_4_update_act) begin
            conv2d_4_dma_flag_1 <= 0;
          end 
          if(conv2d_4_update_act) begin
            conv2d_4_dma_flag_1 <= cparam_conv2d_4_dma_flag_conds_1;
          end 
          if(conv2d_4_update_act && (conv2d_4_row_count >= cparam_conv2d_4_max_row_count)) begin
            conv2d_4_dma_flag_1 <= 1;
          end 
          if(!conv2d_4_update_act) begin
            conv2d_4_dma_flag_2 <= 0;
          end 
          if(conv2d_4_update_act) begin
            conv2d_4_dma_flag_2 <= cparam_conv2d_4_dma_flag_conds_2;
          end 
          if(conv2d_4_update_act && (conv2d_4_row_count >= cparam_conv2d_4_max_row_count)) begin
            conv2d_4_dma_flag_2 <= 1;
          end 
          if(conv2d_4_update_act) begin
            conv2d_4_row_count <= conv2d_4_row_count + cparam_conv2d_4_stride_row_par_row;
          end 
          if(conv2d_4_update_act && (conv2d_4_row_count >= cparam_conv2d_4_max_row_count)) begin
            conv2d_4_row_count <= 0;
            conv2d_4_bat_count <= conv2d_4_bat_count + 1;
          end 
          if(conv2d_4_update_act && (conv2d_4_row_count >= cparam_conv2d_4_max_row_count) && (conv2d_4_bat_count >= cparam_conv2d_4_max_bat_count)) begin
            conv2d_4_bat_count <= 0;
          end 
          if(conv2d_4_update_act && (cparam_conv2d_4_stride_row_par_row < 3)) begin
            conv2d_4_row_select <= conv2d_4_row_select + cparam_conv2d_4_stride_row_par_row;
            conv2d_4_prev_row_select <= conv2d_4_row_select;
          end 
          if(conv2d_4_update_act && (cparam_conv2d_4_stride_row_par_row < 3) && (conv2d_4_row_select + cparam_conv2d_4_stride_row_par_row >= 3)) begin
            conv2d_4_row_select <= conv2d_4_row_select - (3 - cparam_conv2d_4_stride_row_par_row);
            conv2d_4_prev_row_select <= conv2d_4_row_select;
          end 
          if(conv2d_4_update_act && !(cparam_conv2d_4_stride_row_par_row < 3)) begin
            conv2d_4_row_select <= 0;
            conv2d_4_prev_row_select <= 0;
          end 
          if(conv2d_4_update_act && (conv2d_4_row_count >= cparam_conv2d_4_max_row_count)) begin
            conv2d_4_row_select <= 0;
            conv2d_4_prev_row_select <= 0;
          end 
          if(conv2d_4_update_act && conv2d_4_mux_next_dma_flag_0) begin
            conv2d_4_act_page_comp_offset_0 <= conv2d_4_act_page_comp_offset_0 + cparam_conv2d_4_act_read_step;
            conv2d_4_act_page_dma_offset_0 <= conv2d_4_act_page_dma_offset_0 + cparam_conv2d_4_act_read_step;
          end 
          if(conv2d_4_update_act && conv2d_4_mux_next_dma_flag_0 && (conv2d_4_act_page_comp_offset_0 + cparam_conv2d_4_act_read_step + cparam_conv2d_4_act_read_step > 512)) begin
            conv2d_4_act_page_comp_offset_0 <= 0;
            conv2d_4_act_page_dma_offset_0 <= 0;
          end 
          if((cparam_conv2d_4_data_stationary == 0) && (conv2d_4_row_count >= cparam_conv2d_4_max_row_count) && (conv2d_4_bat_count >= cparam_conv2d_4_max_bat_count) && cparam_conv2d_4_keep_input) begin
            conv2d_4_act_page_comp_offset_0 <= 0;
            conv2d_4_act_page_dma_offset_0 <= 0;
          end 
          if(conv2d_4_update_act && conv2d_4_mux_next_dma_flag_1) begin
            conv2d_4_act_page_comp_offset_1 <= conv2d_4_act_page_comp_offset_1 + cparam_conv2d_4_act_read_step;
            conv2d_4_act_page_dma_offset_1 <= conv2d_4_act_page_dma_offset_1 + cparam_conv2d_4_act_read_step;
          end 
          if(conv2d_4_update_act && conv2d_4_mux_next_dma_flag_1 && (conv2d_4_act_page_comp_offset_1 + cparam_conv2d_4_act_read_step + cparam_conv2d_4_act_read_step > 512)) begin
            conv2d_4_act_page_comp_offset_1 <= 0;
            conv2d_4_act_page_dma_offset_1 <= 0;
          end 
          if((cparam_conv2d_4_data_stationary == 0) && (conv2d_4_row_count >= cparam_conv2d_4_max_row_count) && (conv2d_4_bat_count >= cparam_conv2d_4_max_bat_count) && cparam_conv2d_4_keep_input) begin
            conv2d_4_act_page_comp_offset_1 <= 0;
            conv2d_4_act_page_dma_offset_1 <= 0;
          end 
          if(conv2d_4_update_act && conv2d_4_mux_next_dma_flag_2) begin
            conv2d_4_act_page_comp_offset_2 <= conv2d_4_act_page_comp_offset_2 + cparam_conv2d_4_act_read_step;
            conv2d_4_act_page_dma_offset_2 <= conv2d_4_act_page_dma_offset_2 + cparam_conv2d_4_act_read_step;
          end 
          if(conv2d_4_update_act && conv2d_4_mux_next_dma_flag_2 && (conv2d_4_act_page_comp_offset_2 + cparam_conv2d_4_act_read_step + cparam_conv2d_4_act_read_step > 512)) begin
            conv2d_4_act_page_comp_offset_2 <= 0;
            conv2d_4_act_page_dma_offset_2 <= 0;
          end 
          if((cparam_conv2d_4_data_stationary == 0) && (conv2d_4_row_count >= cparam_conv2d_4_max_row_count) && (conv2d_4_bat_count >= cparam_conv2d_4_max_bat_count) && cparam_conv2d_4_keep_input) begin
            conv2d_4_act_page_comp_offset_2 <= 0;
            conv2d_4_act_page_dma_offset_2 <= 0;
          end 
          conv2d_4_next_out_write_size <= (conv2d_4_och_count >= cparam_conv2d_4_max_och_count)? cparam_conv2d_4_out_write_size_res : cparam_conv2d_4_out_write_size;
          if(!conv2d_4_skip_write_out) begin
            conv2d_4_write_count <= 0;
            conv2d_4_out_laddr_offset <= 0;
            conv2d_4_out_ram_select <= 0;
          end 
          if((cparam_conv2d_4_data_stationary == 0) && !conv2d_4_skip_write_out) begin
            conv2d_4_out_base_offset_col <= 0;
            conv2d_4_out_base_offset_row <= conv2d_4_out_base_offset_row + cparam_conv2d_4_out_row_step;
            conv2d_4_out_col_count <= 0;
            conv2d_4_out_row_count <= conv2d_4_out_row_count + 1;
          end 
          if((cparam_conv2d_4_data_stationary == 0) && !conv2d_4_skip_write_out && (conv2d_4_prev_row_count >= cparam_conv2d_4_max_row_count)) begin
            conv2d_4_out_base_offset_row <= 0;
            conv2d_4_out_base_offset_bat <= conv2d_4_out_base_offset_bat + cparam_conv2d_4_out_bat_step;
            conv2d_4_out_row_count <= 0;
          end 
          if((cparam_conv2d_4_data_stationary == 0) && !conv2d_4_skip_write_out && (conv2d_4_prev_row_count >= cparam_conv2d_4_max_row_count) && (conv2d_4_prev_bat_count >= cparam_conv2d_4_max_bat_count)) begin
            conv2d_4_out_base_offset_bat <= 0;
            conv2d_4_out_base_offset_och <= conv2d_4_out_base_offset_och + cparam_conv2d_4_out_och_step;
          end 
          if((cparam_conv2d_4_data_stationary == 1) && (conv2d_4_prev_och_count >= cparam_conv2d_4_max_och_count) && !conv2d_4_skip_write_out) begin
            conv2d_4_out_base_offset_row <= conv2d_4_out_base_offset_row + cparam_conv2d_4_out_row_step;
          end 
          if((cparam_conv2d_4_data_stationary == 0) && !conv2d_4_out_page) begin
            conv2d_4_out_page_comp_offset <= 256;
            conv2d_4_out_page_dma_offset <= 0;
            conv2d_4_out_page <= 1;
          end 
          if((cparam_conv2d_4_data_stationary == 0) && conv2d_4_out_page) begin
            conv2d_4_out_page_comp_offset <= 0;
            conv2d_4_out_page_dma_offset <= 256;
            conv2d_4_out_page <= 0;
          end 
          if((cparam_conv2d_4_data_stationary == 1) && (conv2d_4_och_count >= cparam_conv2d_4_max_och_count) && !conv2d_4_out_page) begin
            conv2d_4_out_page_comp_offset <= 256;
            conv2d_4_out_page_dma_offset <= 0;
            conv2d_4_out_page <= 1;
          end 
          if((cparam_conv2d_4_data_stationary == 1) && (conv2d_4_och_count >= cparam_conv2d_4_max_och_count) && conv2d_4_out_page) begin
            conv2d_4_out_page_comp_offset <= 0;
            conv2d_4_out_page_dma_offset <= 256;
            conv2d_4_out_page <= 0;
          end 
          conv2d_4_prev_row_count <= conv2d_4_row_count;
          conv2d_4_prev_bat_count <= conv2d_4_bat_count;
          conv2d_4_prev_och_count <= conv2d_4_och_count;
          if((conv2d_4_row_count >= cparam_conv2d_4_max_row_count) && (conv2d_4_bat_count >= cparam_conv2d_4_max_bat_count) && (conv2d_4_och_count >= cparam_conv2d_4_max_och_count)) begin
            conv2d_4_skip_read_filter <= 1;
          end 
          if((cparam_conv2d_4_data_stationary == 1) && cparam_conv2d_4_keep_filter) begin
            conv2d_4_skip_read_filter <= 1;
          end 
          if((conv2d_4_row_count >= cparam_conv2d_4_max_row_count) && (conv2d_4_bat_count >= cparam_conv2d_4_max_bat_count) && (conv2d_4_och_count >= cparam_conv2d_4_max_och_count)) begin
            conv2d_4_skip_read_act <= 1;
          end 
          if((cparam_conv2d_4_data_stationary == 0) && (conv2d_4_row_count >= cparam_conv2d_4_max_row_count) && (conv2d_4_bat_count >= cparam_conv2d_4_max_bat_count) && cparam_conv2d_4_keep_input) begin
            conv2d_4_skip_read_act <= 1;
          end 
          if((conv2d_4_row_count >= cparam_conv2d_4_max_row_count) && (conv2d_4_bat_count >= cparam_conv2d_4_max_bat_count) && (conv2d_4_och_count >= cparam_conv2d_4_max_och_count)) begin
            conv2d_4_skip_comp <= 1;
          end 
          if(conv2d_4_skip_write_out && (conv2d_4_prev_row_count == 0) && (conv2d_4_prev_bat_count == 0) && (conv2d_4_prev_och_count == 0)) begin
            conv2d_4_skip_write_out <= 0;
          end 
          if(cparam_conv2d_4_data_stationary == 0) begin
            control_conv2d_4 <= control_conv2d_4_12;
          end 
          if((cparam_conv2d_4_data_stationary == 0) && (conv2d_4_row_count >= cparam_conv2d_4_max_row_count) && (conv2d_4_bat_count >= cparam_conv2d_4_max_bat_count)) begin
            control_conv2d_4 <= control_conv2d_4_7;
          end 
          if(cparam_conv2d_4_data_stationary == 1) begin
            control_conv2d_4 <= control_conv2d_4_7;
          end 
          if((cparam_conv2d_4_data_stationary == 1) && (conv2d_4_och_count >= cparam_conv2d_4_max_och_count)) begin
            control_conv2d_4 <= control_conv2d_4_12;
          end 
          if(!conv2d_4_skip_write_out && (conv2d_4_prev_och_count >= cparam_conv2d_4_max_och_count) && (conv2d_4_prev_row_count >= cparam_conv2d_4_max_row_count) && (conv2d_4_prev_bat_count >= cparam_conv2d_4_max_bat_count)) begin
            control_conv2d_4 <= control_conv2d_4_33;
          end 
        end
        control_conv2d_4_33: begin
          if(_maxi_write_idle && !_maxi_has_outstanding_write) begin
            control_conv2d_4 <= control_conv2d_4_34;
          end 
        end
        control_conv2d_4_34: begin
          if(main_fsm == 13) begin
            _control_conv2d_4_called <= 0;
          end 
          if(main_fsm == 13) begin
            control_conv2d_4 <= control_conv2d_4_init;
          end 
        end
      endcase
    end
  end

  localparam _maxi_read_req_fsm_1 = 1;

  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _maxi_read_req_fsm <= _maxi_read_req_fsm_init;
      _maxi_read_cont <= 0;
    end else begin
      case(_maxi_read_req_fsm)
        _maxi_read_req_fsm_init: begin
          if((_maxi_read_req_fsm == 0) && (_maxi_read_start || _maxi_read_cont) && !_maxi_read_req_fifo_almost_full) begin
            _maxi_read_req_fsm <= _maxi_read_req_fsm_1;
          end 
        end
        _maxi_read_req_fsm_1: begin
          if(maxi_arready || !maxi_arvalid) begin
            _maxi_read_cont <= 1;
          end 
          if((maxi_arready || !maxi_arvalid) && (_maxi_read_global_size == 0)) begin
            _maxi_read_cont <= 0;
          end 
          if(maxi_arready || !maxi_arvalid) begin
            _maxi_read_req_fsm <= _maxi_read_req_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam _maxi_read_data_fsm_1 = 1;
  localparam _maxi_read_data_fsm_2 = 2;

  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
    end else begin
      case(_maxi_read_data_fsm)
        _maxi_read_data_fsm_init: begin
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 2)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 3)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 4)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 5)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 6)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 7)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 8)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 9)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
          if(!_maxi_read_data_busy && !_maxi_read_req_fifo_empty && (_maxi_read_op_sel_fifo == 10)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_1;
          end 
        end
        _maxi_read_data_fsm_1: begin
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
          _maxi_read_data_fsm <= _maxi_read_data_fsm_2;
        end
        _maxi_read_data_fsm_2: begin
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
          if(_maxi_rvalid_sb_0 && (_maxi_read_local_size_buf <= 1)) begin
            _maxi_read_data_fsm <= _maxi_read_data_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_31_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_31 <= write_burst_packed_fsm_31_init;
      write_burst_packed_addr_79 <= 0;
      write_burst_packed_stride_80 <= 0;
      write_burst_packed_length_81 <= 0;
      write_burst_packed_done_82 <= 0;
    end else begin
      case(write_burst_packed_fsm_31)
        write_burst_packed_fsm_31_init: begin
          write_burst_packed_addr_79 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_80 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_81 <= _maxi_read_local_size_buf;
          write_burst_packed_done_82 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 1) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_31 <= write_burst_packed_fsm_31_1;
          end 
        end
        write_burst_packed_fsm_31_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_packed_addr_79 <= write_burst_packed_addr_79 + write_burst_packed_stride_80;
            write_burst_packed_length_81 <= write_burst_packed_length_81 - 1;
            write_burst_packed_done_82 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_packed_length_81 <= 1)) begin
            write_burst_packed_done_82 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_packed_done_82 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_packed_length_81 <= 1)) begin
            write_burst_packed_fsm_31 <= write_burst_packed_fsm_31_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_packed_fsm_31 <= write_burst_packed_fsm_31_init;
          end 
          if(0) begin
            write_burst_packed_fsm_31 <= write_burst_packed_fsm_31_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_32_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_32 <= write_burst_packed_fsm_32_init;
      write_burst_packed_addr_92 <= 0;
      write_burst_packed_stride_93 <= 0;
      write_burst_packed_length_94 <= 0;
      write_burst_packed_done_95 <= 0;
    end else begin
      case(write_burst_packed_fsm_32)
        write_burst_packed_fsm_32_init: begin
          write_burst_packed_addr_92 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_93 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_94 <= _maxi_read_local_size_buf;
          write_burst_packed_done_95 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 2) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_32 <= write_burst_packed_fsm_32_1;
          end 
        end
        write_burst_packed_fsm_32_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_packed_addr_92 <= write_burst_packed_addr_92 + write_burst_packed_stride_93;
            write_burst_packed_length_94 <= write_burst_packed_length_94 - 1;
            write_burst_packed_done_95 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_packed_length_94 <= 1)) begin
            write_burst_packed_done_95 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_packed_done_95 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_packed_length_94 <= 1)) begin
            write_burst_packed_fsm_32 <= write_burst_packed_fsm_32_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_packed_fsm_32 <= write_burst_packed_fsm_32_init;
          end 
          if(0) begin
            write_burst_packed_fsm_32 <= write_burst_packed_fsm_32_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_33_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_33 <= write_burst_packed_fsm_33_init;
      write_burst_packed_addr_110 <= 0;
      write_burst_packed_stride_111 <= 0;
      write_burst_packed_length_112 <= 0;
      write_burst_packed_done_113 <= 0;
    end else begin
      case(write_burst_packed_fsm_33)
        write_burst_packed_fsm_33_init: begin
          write_burst_packed_addr_110 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_111 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_112 <= _maxi_read_local_size_buf;
          write_burst_packed_done_113 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_33 <= write_burst_packed_fsm_33_1;
          end 
        end
        write_burst_packed_fsm_33_1: begin
          if(write_burst_block_ram_wvalid_108) begin
            write_burst_packed_addr_110 <= write_burst_packed_addr_110 + write_burst_packed_stride_111;
            write_burst_packed_length_112 <= write_burst_packed_length_112 - 1;
            write_burst_packed_done_113 <= 0;
          end 
          if(write_burst_block_ram_wvalid_108 && (write_burst_packed_length_112 <= 1)) begin
            write_burst_packed_done_113 <= 1;
          end 
          if(write_burst_block_ram_wvalid_108 && 0) begin
            write_burst_packed_done_113 <= 1;
          end 
          if(write_burst_block_ram_wvalid_108 && (write_burst_packed_length_112 <= 1)) begin
            write_burst_packed_fsm_33 <= write_burst_packed_fsm_33_init;
          end 
          if(write_burst_block_ram_wvalid_108 && 0) begin
            write_burst_packed_fsm_33 <= write_burst_packed_fsm_33_init;
          end 
          if(write_burst_block_ram_wquit_109) begin
            write_burst_packed_fsm_33 <= write_burst_packed_fsm_33_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_34_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_34 <= write_burst_packed_fsm_34_init;
      write_burst_packed_addr_120 <= 0;
      write_burst_packed_stride_121 <= 0;
      write_burst_packed_length_122 <= 0;
      write_burst_packed_done_123 <= 0;
    end else begin
      case(write_burst_packed_fsm_34)
        write_burst_packed_fsm_34_init: begin
          write_burst_packed_addr_120 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_121 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_122 <= _maxi_read_local_size_buf;
          write_burst_packed_done_123 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_34 <= write_burst_packed_fsm_34_1;
          end 
        end
        write_burst_packed_fsm_34_1: begin
          if(write_burst_block_ram_wvalid_118) begin
            write_burst_packed_addr_120 <= write_burst_packed_addr_120 + write_burst_packed_stride_121;
            write_burst_packed_length_122 <= write_burst_packed_length_122 - 1;
            write_burst_packed_done_123 <= 0;
          end 
          if(write_burst_block_ram_wvalid_118 && (write_burst_packed_length_122 <= 1)) begin
            write_burst_packed_done_123 <= 1;
          end 
          if(write_burst_block_ram_wvalid_118 && 0) begin
            write_burst_packed_done_123 <= 1;
          end 
          if(write_burst_block_ram_wvalid_118 && (write_burst_packed_length_122 <= 1)) begin
            write_burst_packed_fsm_34 <= write_burst_packed_fsm_34_init;
          end 
          if(write_burst_block_ram_wvalid_118 && 0) begin
            write_burst_packed_fsm_34 <= write_burst_packed_fsm_34_init;
          end 
          if(write_burst_block_ram_wquit_119) begin
            write_burst_packed_fsm_34 <= write_burst_packed_fsm_34_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_35_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_35 <= write_burst_packed_fsm_35_init;
      write_burst_packed_addr_130 <= 0;
      write_burst_packed_stride_131 <= 0;
      write_burst_packed_length_132 <= 0;
      write_burst_packed_done_133 <= 0;
    end else begin
      case(write_burst_packed_fsm_35)
        write_burst_packed_fsm_35_init: begin
          write_burst_packed_addr_130 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_131 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_132 <= _maxi_read_local_size_buf;
          write_burst_packed_done_133 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_35 <= write_burst_packed_fsm_35_1;
          end 
        end
        write_burst_packed_fsm_35_1: begin
          if(write_burst_block_ram_wvalid_128) begin
            write_burst_packed_addr_130 <= write_burst_packed_addr_130 + write_burst_packed_stride_131;
            write_burst_packed_length_132 <= write_burst_packed_length_132 - 1;
            write_burst_packed_done_133 <= 0;
          end 
          if(write_burst_block_ram_wvalid_128 && (write_burst_packed_length_132 <= 1)) begin
            write_burst_packed_done_133 <= 1;
          end 
          if(write_burst_block_ram_wvalid_128 && 0) begin
            write_burst_packed_done_133 <= 1;
          end 
          if(write_burst_block_ram_wvalid_128 && (write_burst_packed_length_132 <= 1)) begin
            write_burst_packed_fsm_35 <= write_burst_packed_fsm_35_init;
          end 
          if(write_burst_block_ram_wvalid_128 && 0) begin
            write_burst_packed_fsm_35 <= write_burst_packed_fsm_35_init;
          end 
          if(write_burst_block_ram_wquit_129) begin
            write_burst_packed_fsm_35 <= write_burst_packed_fsm_35_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_36_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_36 <= write_burst_packed_fsm_36_init;
      write_burst_packed_addr_140 <= 0;
      write_burst_packed_stride_141 <= 0;
      write_burst_packed_length_142 <= 0;
      write_burst_packed_done_143 <= 0;
    end else begin
      case(write_burst_packed_fsm_36)
        write_burst_packed_fsm_36_init: begin
          write_burst_packed_addr_140 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_141 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_142 <= _maxi_read_local_size_buf;
          write_burst_packed_done_143 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_36 <= write_burst_packed_fsm_36_1;
          end 
        end
        write_burst_packed_fsm_36_1: begin
          if(write_burst_block_ram_wvalid_138) begin
            write_burst_packed_addr_140 <= write_burst_packed_addr_140 + write_burst_packed_stride_141;
            write_burst_packed_length_142 <= write_burst_packed_length_142 - 1;
            write_burst_packed_done_143 <= 0;
          end 
          if(write_burst_block_ram_wvalid_138 && (write_burst_packed_length_142 <= 1)) begin
            write_burst_packed_done_143 <= 1;
          end 
          if(write_burst_block_ram_wvalid_138 && 0) begin
            write_burst_packed_done_143 <= 1;
          end 
          if(write_burst_block_ram_wvalid_138 && (write_burst_packed_length_142 <= 1)) begin
            write_burst_packed_fsm_36 <= write_burst_packed_fsm_36_init;
          end 
          if(write_burst_block_ram_wvalid_138 && 0) begin
            write_burst_packed_fsm_36 <= write_burst_packed_fsm_36_init;
          end 
          if(write_burst_block_ram_wquit_139) begin
            write_burst_packed_fsm_36 <= write_burst_packed_fsm_36_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_37_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_37 <= write_burst_packed_fsm_37_init;
      write_burst_packed_addr_150 <= 0;
      write_burst_packed_stride_151 <= 0;
      write_burst_packed_length_152 <= 0;
      write_burst_packed_done_153 <= 0;
    end else begin
      case(write_burst_packed_fsm_37)
        write_burst_packed_fsm_37_init: begin
          write_burst_packed_addr_150 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_151 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_152 <= _maxi_read_local_size_buf;
          write_burst_packed_done_153 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_37 <= write_burst_packed_fsm_37_1;
          end 
        end
        write_burst_packed_fsm_37_1: begin
          if(write_burst_block_ram_wvalid_148) begin
            write_burst_packed_addr_150 <= write_burst_packed_addr_150 + write_burst_packed_stride_151;
            write_burst_packed_length_152 <= write_burst_packed_length_152 - 1;
            write_burst_packed_done_153 <= 0;
          end 
          if(write_burst_block_ram_wvalid_148 && (write_burst_packed_length_152 <= 1)) begin
            write_burst_packed_done_153 <= 1;
          end 
          if(write_burst_block_ram_wvalid_148 && 0) begin
            write_burst_packed_done_153 <= 1;
          end 
          if(write_burst_block_ram_wvalid_148 && (write_burst_packed_length_152 <= 1)) begin
            write_burst_packed_fsm_37 <= write_burst_packed_fsm_37_init;
          end 
          if(write_burst_block_ram_wvalid_148 && 0) begin
            write_burst_packed_fsm_37 <= write_burst_packed_fsm_37_init;
          end 
          if(write_burst_block_ram_wquit_149) begin
            write_burst_packed_fsm_37 <= write_burst_packed_fsm_37_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_38_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_38 <= write_burst_packed_fsm_38_init;
      write_burst_packed_addr_160 <= 0;
      write_burst_packed_stride_161 <= 0;
      write_burst_packed_length_162 <= 0;
      write_burst_packed_done_163 <= 0;
    end else begin
      case(write_burst_packed_fsm_38)
        write_burst_packed_fsm_38_init: begin
          write_burst_packed_addr_160 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_161 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_162 <= _maxi_read_local_size_buf;
          write_burst_packed_done_163 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_38 <= write_burst_packed_fsm_38_1;
          end 
        end
        write_burst_packed_fsm_38_1: begin
          if(write_burst_block_ram_wvalid_158) begin
            write_burst_packed_addr_160 <= write_burst_packed_addr_160 + write_burst_packed_stride_161;
            write_burst_packed_length_162 <= write_burst_packed_length_162 - 1;
            write_burst_packed_done_163 <= 0;
          end 
          if(write_burst_block_ram_wvalid_158 && (write_burst_packed_length_162 <= 1)) begin
            write_burst_packed_done_163 <= 1;
          end 
          if(write_burst_block_ram_wvalid_158 && 0) begin
            write_burst_packed_done_163 <= 1;
          end 
          if(write_burst_block_ram_wvalid_158 && (write_burst_packed_length_162 <= 1)) begin
            write_burst_packed_fsm_38 <= write_burst_packed_fsm_38_init;
          end 
          if(write_burst_block_ram_wvalid_158 && 0) begin
            write_burst_packed_fsm_38 <= write_burst_packed_fsm_38_init;
          end 
          if(write_burst_block_ram_wquit_159) begin
            write_burst_packed_fsm_38 <= write_burst_packed_fsm_38_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_39_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_39 <= write_burst_packed_fsm_39_init;
      write_burst_packed_addr_170 <= 0;
      write_burst_packed_stride_171 <= 0;
      write_burst_packed_length_172 <= 0;
      write_burst_packed_done_173 <= 0;
    end else begin
      case(write_burst_packed_fsm_39)
        write_burst_packed_fsm_39_init: begin
          write_burst_packed_addr_170 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_171 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_172 <= _maxi_read_local_size_buf;
          write_burst_packed_done_173 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_39 <= write_burst_packed_fsm_39_1;
          end 
        end
        write_burst_packed_fsm_39_1: begin
          if(write_burst_block_ram_wvalid_168) begin
            write_burst_packed_addr_170 <= write_burst_packed_addr_170 + write_burst_packed_stride_171;
            write_burst_packed_length_172 <= write_burst_packed_length_172 - 1;
            write_burst_packed_done_173 <= 0;
          end 
          if(write_burst_block_ram_wvalid_168 && (write_burst_packed_length_172 <= 1)) begin
            write_burst_packed_done_173 <= 1;
          end 
          if(write_burst_block_ram_wvalid_168 && 0) begin
            write_burst_packed_done_173 <= 1;
          end 
          if(write_burst_block_ram_wvalid_168 && (write_burst_packed_length_172 <= 1)) begin
            write_burst_packed_fsm_39 <= write_burst_packed_fsm_39_init;
          end 
          if(write_burst_block_ram_wvalid_168 && 0) begin
            write_burst_packed_fsm_39 <= write_burst_packed_fsm_39_init;
          end 
          if(write_burst_block_ram_wquit_169) begin
            write_burst_packed_fsm_39 <= write_burst_packed_fsm_39_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_40_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_40 <= write_burst_packed_fsm_40_init;
      write_burst_packed_addr_180 <= 0;
      write_burst_packed_stride_181 <= 0;
      write_burst_packed_length_182 <= 0;
      write_burst_packed_done_183 <= 0;
    end else begin
      case(write_burst_packed_fsm_40)
        write_burst_packed_fsm_40_init: begin
          write_burst_packed_addr_180 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_181 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_182 <= _maxi_read_local_size_buf;
          write_burst_packed_done_183 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_40 <= write_burst_packed_fsm_40_1;
          end 
        end
        write_burst_packed_fsm_40_1: begin
          if(write_burst_block_ram_wvalid_178) begin
            write_burst_packed_addr_180 <= write_burst_packed_addr_180 + write_burst_packed_stride_181;
            write_burst_packed_length_182 <= write_burst_packed_length_182 - 1;
            write_burst_packed_done_183 <= 0;
          end 
          if(write_burst_block_ram_wvalid_178 && (write_burst_packed_length_182 <= 1)) begin
            write_burst_packed_done_183 <= 1;
          end 
          if(write_burst_block_ram_wvalid_178 && 0) begin
            write_burst_packed_done_183 <= 1;
          end 
          if(write_burst_block_ram_wvalid_178 && (write_burst_packed_length_182 <= 1)) begin
            write_burst_packed_fsm_40 <= write_burst_packed_fsm_40_init;
          end 
          if(write_burst_block_ram_wvalid_178 && 0) begin
            write_burst_packed_fsm_40 <= write_burst_packed_fsm_40_init;
          end 
          if(write_burst_block_ram_wquit_179) begin
            write_burst_packed_fsm_40 <= write_burst_packed_fsm_40_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_41_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_41 <= write_burst_packed_fsm_41_init;
      write_burst_packed_addr_190 <= 0;
      write_burst_packed_stride_191 <= 0;
      write_burst_packed_length_192 <= 0;
      write_burst_packed_done_193 <= 0;
    end else begin
      case(write_burst_packed_fsm_41)
        write_burst_packed_fsm_41_init: begin
          write_burst_packed_addr_190 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_191 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_192 <= _maxi_read_local_size_buf;
          write_burst_packed_done_193 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_41 <= write_burst_packed_fsm_41_1;
          end 
        end
        write_burst_packed_fsm_41_1: begin
          if(write_burst_block_ram_wvalid_188) begin
            write_burst_packed_addr_190 <= write_burst_packed_addr_190 + write_burst_packed_stride_191;
            write_burst_packed_length_192 <= write_burst_packed_length_192 - 1;
            write_burst_packed_done_193 <= 0;
          end 
          if(write_burst_block_ram_wvalid_188 && (write_burst_packed_length_192 <= 1)) begin
            write_burst_packed_done_193 <= 1;
          end 
          if(write_burst_block_ram_wvalid_188 && 0) begin
            write_burst_packed_done_193 <= 1;
          end 
          if(write_burst_block_ram_wvalid_188 && (write_burst_packed_length_192 <= 1)) begin
            write_burst_packed_fsm_41 <= write_burst_packed_fsm_41_init;
          end 
          if(write_burst_block_ram_wvalid_188 && 0) begin
            write_burst_packed_fsm_41 <= write_burst_packed_fsm_41_init;
          end 
          if(write_burst_block_ram_wquit_189) begin
            write_burst_packed_fsm_41 <= write_burst_packed_fsm_41_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_block_fsm_42_1 = 1;
  localparam write_burst_block_fsm_42_2 = 2;
  localparam write_burst_block_fsm_42_3 = 3;
  localparam write_burst_block_fsm_42_4 = 4;
  localparam write_burst_block_fsm_42_5 = 5;
  localparam write_burst_block_fsm_42_6 = 6;
  localparam write_burst_block_fsm_42_7 = 7;
  localparam write_burst_block_fsm_42_8 = 8;
  localparam write_burst_block_fsm_42_9 = 9;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_block_fsm_42 <= write_burst_block_fsm_42_init;
      write_burst_block_length_198 <= 0;
      write_burst_block_blocksize_199 <= 0;
      write_burst_block_done_200 <= 0;
      write_burst_block_count_201 <= 0;
    end else begin
      case(write_burst_block_fsm_42)
        write_burst_block_fsm_42_init: begin
          write_burst_block_length_198 <= _maxi_read_local_size_buf;
          write_burst_block_blocksize_199 <= _maxi_read_local_blocksize_buf;
          write_burst_block_done_200 <= 0;
          write_burst_block_count_201 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 3) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_block_fsm_42 <= write_burst_block_fsm_42_1;
          end 
        end
        write_burst_block_fsm_42_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_198 <= write_burst_block_length_198 - 1;
            write_burst_block_done_200 <= 0;
            write_burst_block_count_201 <= write_burst_block_count_201 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1)) begin
            write_burst_block_done_200 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_200 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_201 == write_burst_block_blocksize_199 - 1)) begin
            write_burst_block_count_201 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_201 == write_burst_block_blocksize_199 - 1)) begin
            write_burst_block_fsm_42 <= write_burst_block_fsm_42_2;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1)) begin
            write_burst_block_fsm_42 <= write_burst_block_fsm_42_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_42 <= write_burst_block_fsm_42_init;
          end 
          if(0) begin
            write_burst_block_fsm_42 <= write_burst_block_fsm_42_init;
          end 
        end
        write_burst_block_fsm_42_2: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_198 <= write_burst_block_length_198 - 1;
            write_burst_block_done_200 <= 0;
            write_burst_block_count_201 <= write_burst_block_count_201 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1)) begin
            write_burst_block_done_200 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_200 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_201 == write_burst_block_blocksize_199 - 1)) begin
            write_burst_block_count_201 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_201 == write_burst_block_blocksize_199 - 1)) begin
            write_burst_block_fsm_42 <= write_burst_block_fsm_42_3;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1)) begin
            write_burst_block_fsm_42 <= write_burst_block_fsm_42_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_42 <= write_burst_block_fsm_42_init;
          end 
          if(0) begin
            write_burst_block_fsm_42 <= write_burst_block_fsm_42_init;
          end 
        end
        write_burst_block_fsm_42_3: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_198 <= write_burst_block_length_198 - 1;
            write_burst_block_done_200 <= 0;
            write_burst_block_count_201 <= write_burst_block_count_201 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1)) begin
            write_burst_block_done_200 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_200 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_201 == write_burst_block_blocksize_199 - 1)) begin
            write_burst_block_count_201 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_201 == write_burst_block_blocksize_199 - 1)) begin
            write_burst_block_fsm_42 <= write_burst_block_fsm_42_4;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1)) begin
            write_burst_block_fsm_42 <= write_burst_block_fsm_42_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_42 <= write_burst_block_fsm_42_init;
          end 
          if(0) begin
            write_burst_block_fsm_42 <= write_burst_block_fsm_42_init;
          end 
        end
        write_burst_block_fsm_42_4: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_198 <= write_burst_block_length_198 - 1;
            write_burst_block_done_200 <= 0;
            write_burst_block_count_201 <= write_burst_block_count_201 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1)) begin
            write_burst_block_done_200 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_200 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_201 == write_burst_block_blocksize_199 - 1)) begin
            write_burst_block_count_201 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_201 == write_burst_block_blocksize_199 - 1)) begin
            write_burst_block_fsm_42 <= write_burst_block_fsm_42_5;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1)) begin
            write_burst_block_fsm_42 <= write_burst_block_fsm_42_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_42 <= write_burst_block_fsm_42_init;
          end 
          if(0) begin
            write_burst_block_fsm_42 <= write_burst_block_fsm_42_init;
          end 
        end
        write_burst_block_fsm_42_5: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_198 <= write_burst_block_length_198 - 1;
            write_burst_block_done_200 <= 0;
            write_burst_block_count_201 <= write_burst_block_count_201 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1)) begin
            write_burst_block_done_200 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_200 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_201 == write_burst_block_blocksize_199 - 1)) begin
            write_burst_block_count_201 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_201 == write_burst_block_blocksize_199 - 1)) begin
            write_burst_block_fsm_42 <= write_burst_block_fsm_42_6;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1)) begin
            write_burst_block_fsm_42 <= write_burst_block_fsm_42_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_42 <= write_burst_block_fsm_42_init;
          end 
          if(0) begin
            write_burst_block_fsm_42 <= write_burst_block_fsm_42_init;
          end 
        end
        write_burst_block_fsm_42_6: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_198 <= write_burst_block_length_198 - 1;
            write_burst_block_done_200 <= 0;
            write_burst_block_count_201 <= write_burst_block_count_201 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1)) begin
            write_burst_block_done_200 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_200 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_201 == write_burst_block_blocksize_199 - 1)) begin
            write_burst_block_count_201 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_201 == write_burst_block_blocksize_199 - 1)) begin
            write_burst_block_fsm_42 <= write_burst_block_fsm_42_7;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1)) begin
            write_burst_block_fsm_42 <= write_burst_block_fsm_42_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_42 <= write_burst_block_fsm_42_init;
          end 
          if(0) begin
            write_burst_block_fsm_42 <= write_burst_block_fsm_42_init;
          end 
        end
        write_burst_block_fsm_42_7: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_198 <= write_burst_block_length_198 - 1;
            write_burst_block_done_200 <= 0;
            write_burst_block_count_201 <= write_burst_block_count_201 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1)) begin
            write_burst_block_done_200 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_200 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_201 == write_burst_block_blocksize_199 - 1)) begin
            write_burst_block_count_201 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_201 == write_burst_block_blocksize_199 - 1)) begin
            write_burst_block_fsm_42 <= write_burst_block_fsm_42_8;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1)) begin
            write_burst_block_fsm_42 <= write_burst_block_fsm_42_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_42 <= write_burst_block_fsm_42_init;
          end 
          if(0) begin
            write_burst_block_fsm_42 <= write_burst_block_fsm_42_init;
          end 
        end
        write_burst_block_fsm_42_8: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_198 <= write_burst_block_length_198 - 1;
            write_burst_block_done_200 <= 0;
            write_burst_block_count_201 <= write_burst_block_count_201 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1)) begin
            write_burst_block_done_200 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_200 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_201 == write_burst_block_blocksize_199 - 1)) begin
            write_burst_block_count_201 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_201 == write_burst_block_blocksize_199 - 1)) begin
            write_burst_block_fsm_42 <= write_burst_block_fsm_42_9;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1)) begin
            write_burst_block_fsm_42 <= write_burst_block_fsm_42_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_42 <= write_burst_block_fsm_42_init;
          end 
          if(0) begin
            write_burst_block_fsm_42 <= write_burst_block_fsm_42_init;
          end 
        end
        write_burst_block_fsm_42_9: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_198 <= write_burst_block_length_198 - 1;
            write_burst_block_done_200 <= 0;
            write_burst_block_count_201 <= write_burst_block_count_201 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1)) begin
            write_burst_block_done_200 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_200 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_201 == write_burst_block_blocksize_199 - 1)) begin
            write_burst_block_count_201 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_201 == write_burst_block_blocksize_199 - 1)) begin
            write_burst_block_fsm_42 <= write_burst_block_fsm_42_1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_198 <= 1)) begin
            write_burst_block_fsm_42 <= write_burst_block_fsm_42_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_42 <= write_burst_block_fsm_42_init;
          end 
          if(0) begin
            write_burst_block_fsm_42 <= write_burst_block_fsm_42_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_43_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_43 <= write_burst_packed_fsm_43_init;
      write_burst_packed_addr_212 <= 0;
      write_burst_packed_stride_213 <= 0;
      write_burst_packed_length_214 <= 0;
      write_burst_packed_done_215 <= 0;
    end else begin
      case(write_burst_packed_fsm_43)
        write_burst_packed_fsm_43_init: begin
          write_burst_packed_addr_212 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_213 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_214 <= _maxi_read_local_size_buf;
          write_burst_packed_done_215 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 4) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_43 <= write_burst_packed_fsm_43_1;
          end 
        end
        write_burst_packed_fsm_43_1: begin
          if(write_burst_block_ram_wvalid_210) begin
            write_burst_packed_addr_212 <= write_burst_packed_addr_212 + write_burst_packed_stride_213;
            write_burst_packed_length_214 <= write_burst_packed_length_214 - 1;
            write_burst_packed_done_215 <= 0;
          end 
          if(write_burst_block_ram_wvalid_210 && (write_burst_packed_length_214 <= 1)) begin
            write_burst_packed_done_215 <= 1;
          end 
          if(write_burst_block_ram_wvalid_210 && 0) begin
            write_burst_packed_done_215 <= 1;
          end 
          if(write_burst_block_ram_wvalid_210 && (write_burst_packed_length_214 <= 1)) begin
            write_burst_packed_fsm_43 <= write_burst_packed_fsm_43_init;
          end 
          if(write_burst_block_ram_wvalid_210 && 0) begin
            write_burst_packed_fsm_43 <= write_burst_packed_fsm_43_init;
          end 
          if(write_burst_block_ram_wquit_211) begin
            write_burst_packed_fsm_43 <= write_burst_packed_fsm_43_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_44_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_44 <= write_burst_packed_fsm_44_init;
      write_burst_packed_addr_222 <= 0;
      write_burst_packed_stride_223 <= 0;
      write_burst_packed_length_224 <= 0;
      write_burst_packed_done_225 <= 0;
    end else begin
      case(write_burst_packed_fsm_44)
        write_burst_packed_fsm_44_init: begin
          write_burst_packed_addr_222 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_223 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_224 <= _maxi_read_local_size_buf;
          write_burst_packed_done_225 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 4) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_44 <= write_burst_packed_fsm_44_1;
          end 
        end
        write_burst_packed_fsm_44_1: begin
          if(write_burst_block_ram_wvalid_220) begin
            write_burst_packed_addr_222 <= write_burst_packed_addr_222 + write_burst_packed_stride_223;
            write_burst_packed_length_224 <= write_burst_packed_length_224 - 1;
            write_burst_packed_done_225 <= 0;
          end 
          if(write_burst_block_ram_wvalid_220 && (write_burst_packed_length_224 <= 1)) begin
            write_burst_packed_done_225 <= 1;
          end 
          if(write_burst_block_ram_wvalid_220 && 0) begin
            write_burst_packed_done_225 <= 1;
          end 
          if(write_burst_block_ram_wvalid_220 && (write_burst_packed_length_224 <= 1)) begin
            write_burst_packed_fsm_44 <= write_burst_packed_fsm_44_init;
          end 
          if(write_burst_block_ram_wvalid_220 && 0) begin
            write_burst_packed_fsm_44 <= write_burst_packed_fsm_44_init;
          end 
          if(write_burst_block_ram_wquit_221) begin
            write_burst_packed_fsm_44 <= write_burst_packed_fsm_44_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_45_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_45 <= write_burst_packed_fsm_45_init;
      write_burst_packed_addr_232 <= 0;
      write_burst_packed_stride_233 <= 0;
      write_burst_packed_length_234 <= 0;
      write_burst_packed_done_235 <= 0;
    end else begin
      case(write_burst_packed_fsm_45)
        write_burst_packed_fsm_45_init: begin
          write_burst_packed_addr_232 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_233 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_234 <= _maxi_read_local_size_buf;
          write_burst_packed_done_235 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 4) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_45 <= write_burst_packed_fsm_45_1;
          end 
        end
        write_burst_packed_fsm_45_1: begin
          if(write_burst_block_ram_wvalid_230) begin
            write_burst_packed_addr_232 <= write_burst_packed_addr_232 + write_burst_packed_stride_233;
            write_burst_packed_length_234 <= write_burst_packed_length_234 - 1;
            write_burst_packed_done_235 <= 0;
          end 
          if(write_burst_block_ram_wvalid_230 && (write_burst_packed_length_234 <= 1)) begin
            write_burst_packed_done_235 <= 1;
          end 
          if(write_burst_block_ram_wvalid_230 && 0) begin
            write_burst_packed_done_235 <= 1;
          end 
          if(write_burst_block_ram_wvalid_230 && (write_burst_packed_length_234 <= 1)) begin
            write_burst_packed_fsm_45 <= write_burst_packed_fsm_45_init;
          end 
          if(write_burst_block_ram_wvalid_230 && 0) begin
            write_burst_packed_fsm_45 <= write_burst_packed_fsm_45_init;
          end 
          if(write_burst_block_ram_wquit_231) begin
            write_burst_packed_fsm_45 <= write_burst_packed_fsm_45_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_block_fsm_46_1 = 1;
  localparam write_burst_block_fsm_46_2 = 2;
  localparam write_burst_block_fsm_46_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_block_fsm_46 <= write_burst_block_fsm_46_init;
      write_burst_block_length_240 <= 0;
      write_burst_block_blocksize_241 <= 0;
      write_burst_block_done_242 <= 0;
      write_burst_block_count_243 <= 0;
    end else begin
      case(write_burst_block_fsm_46)
        write_burst_block_fsm_46_init: begin
          write_burst_block_length_240 <= _maxi_read_local_size_buf;
          write_burst_block_blocksize_241 <= _maxi_read_local_blocksize_buf;
          write_burst_block_done_242 <= 0;
          write_burst_block_count_243 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 4) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_block_fsm_46 <= write_burst_block_fsm_46_1;
          end 
        end
        write_burst_block_fsm_46_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_240 <= write_burst_block_length_240 - 1;
            write_burst_block_done_242 <= 0;
            write_burst_block_count_243 <= write_burst_block_count_243 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_240 <= 1)) begin
            write_burst_block_done_242 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_242 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_243 == write_burst_block_blocksize_241 - 1)) begin
            write_burst_block_count_243 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_243 == write_burst_block_blocksize_241 - 1)) begin
            write_burst_block_fsm_46 <= write_burst_block_fsm_46_2;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_240 <= 1)) begin
            write_burst_block_fsm_46 <= write_burst_block_fsm_46_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_46 <= write_burst_block_fsm_46_init;
          end 
          if(0) begin
            write_burst_block_fsm_46 <= write_burst_block_fsm_46_init;
          end 
        end
        write_burst_block_fsm_46_2: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_240 <= write_burst_block_length_240 - 1;
            write_burst_block_done_242 <= 0;
            write_burst_block_count_243 <= write_burst_block_count_243 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_240 <= 1)) begin
            write_burst_block_done_242 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_242 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_243 == write_burst_block_blocksize_241 - 1)) begin
            write_burst_block_count_243 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_243 == write_burst_block_blocksize_241 - 1)) begin
            write_burst_block_fsm_46 <= write_burst_block_fsm_46_3;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_240 <= 1)) begin
            write_burst_block_fsm_46 <= write_burst_block_fsm_46_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_46 <= write_burst_block_fsm_46_init;
          end 
          if(0) begin
            write_burst_block_fsm_46 <= write_burst_block_fsm_46_init;
          end 
        end
        write_burst_block_fsm_46_3: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_240 <= write_burst_block_length_240 - 1;
            write_burst_block_done_242 <= 0;
            write_burst_block_count_243 <= write_burst_block_count_243 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_240 <= 1)) begin
            write_burst_block_done_242 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_242 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_243 == write_burst_block_blocksize_241 - 1)) begin
            write_burst_block_count_243 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_243 == write_burst_block_blocksize_241 - 1)) begin
            write_burst_block_fsm_46 <= write_burst_block_fsm_46_1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_240 <= 1)) begin
            write_burst_block_fsm_46 <= write_burst_block_fsm_46_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_46 <= write_burst_block_fsm_46_init;
          end 
          if(0) begin
            write_burst_block_fsm_46 <= write_burst_block_fsm_46_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_47_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_47 <= write_burst_packed_fsm_47_init;
      write_burst_packed_addr_254 <= 0;
      write_burst_packed_stride_255 <= 0;
      write_burst_packed_length_256 <= 0;
      write_burst_packed_done_257 <= 0;
    end else begin
      case(write_burst_packed_fsm_47)
        write_burst_packed_fsm_47_init: begin
          write_burst_packed_addr_254 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_255 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_256 <= _maxi_read_local_size_buf;
          write_burst_packed_done_257 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 5) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_47 <= write_burst_packed_fsm_47_1;
          end 
        end
        write_burst_packed_fsm_47_1: begin
          if(write_burst_block_ram_wvalid_252) begin
            write_burst_packed_addr_254 <= write_burst_packed_addr_254 + write_burst_packed_stride_255;
            write_burst_packed_length_256 <= write_burst_packed_length_256 - 1;
            write_burst_packed_done_257 <= 0;
          end 
          if(write_burst_block_ram_wvalid_252 && (write_burst_packed_length_256 <= 1)) begin
            write_burst_packed_done_257 <= 1;
          end 
          if(write_burst_block_ram_wvalid_252 && 0) begin
            write_burst_packed_done_257 <= 1;
          end 
          if(write_burst_block_ram_wvalid_252 && (write_burst_packed_length_256 <= 1)) begin
            write_burst_packed_fsm_47 <= write_burst_packed_fsm_47_init;
          end 
          if(write_burst_block_ram_wvalid_252 && 0) begin
            write_burst_packed_fsm_47 <= write_burst_packed_fsm_47_init;
          end 
          if(write_burst_block_ram_wquit_253) begin
            write_burst_packed_fsm_47 <= write_burst_packed_fsm_47_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_48_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_48 <= write_burst_packed_fsm_48_init;
      write_burst_packed_addr_264 <= 0;
      write_burst_packed_stride_265 <= 0;
      write_burst_packed_length_266 <= 0;
      write_burst_packed_done_267 <= 0;
    end else begin
      case(write_burst_packed_fsm_48)
        write_burst_packed_fsm_48_init: begin
          write_burst_packed_addr_264 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_265 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_266 <= _maxi_read_local_size_buf;
          write_burst_packed_done_267 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 5) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_48 <= write_burst_packed_fsm_48_1;
          end 
        end
        write_burst_packed_fsm_48_1: begin
          if(write_burst_block_ram_wvalid_262) begin
            write_burst_packed_addr_264 <= write_burst_packed_addr_264 + write_burst_packed_stride_265;
            write_burst_packed_length_266 <= write_burst_packed_length_266 - 1;
            write_burst_packed_done_267 <= 0;
          end 
          if(write_burst_block_ram_wvalid_262 && (write_burst_packed_length_266 <= 1)) begin
            write_burst_packed_done_267 <= 1;
          end 
          if(write_burst_block_ram_wvalid_262 && 0) begin
            write_burst_packed_done_267 <= 1;
          end 
          if(write_burst_block_ram_wvalid_262 && (write_burst_packed_length_266 <= 1)) begin
            write_burst_packed_fsm_48 <= write_burst_packed_fsm_48_init;
          end 
          if(write_burst_block_ram_wvalid_262 && 0) begin
            write_burst_packed_fsm_48 <= write_burst_packed_fsm_48_init;
          end 
          if(write_burst_block_ram_wquit_263) begin
            write_burst_packed_fsm_48 <= write_burst_packed_fsm_48_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_49_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_49 <= write_burst_packed_fsm_49_init;
      write_burst_packed_addr_274 <= 0;
      write_burst_packed_stride_275 <= 0;
      write_burst_packed_length_276 <= 0;
      write_burst_packed_done_277 <= 0;
    end else begin
      case(write_burst_packed_fsm_49)
        write_burst_packed_fsm_49_init: begin
          write_burst_packed_addr_274 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_275 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_276 <= _maxi_read_local_size_buf;
          write_burst_packed_done_277 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 5) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_49 <= write_burst_packed_fsm_49_1;
          end 
        end
        write_burst_packed_fsm_49_1: begin
          if(write_burst_block_ram_wvalid_272) begin
            write_burst_packed_addr_274 <= write_burst_packed_addr_274 + write_burst_packed_stride_275;
            write_burst_packed_length_276 <= write_burst_packed_length_276 - 1;
            write_burst_packed_done_277 <= 0;
          end 
          if(write_burst_block_ram_wvalid_272 && (write_burst_packed_length_276 <= 1)) begin
            write_burst_packed_done_277 <= 1;
          end 
          if(write_burst_block_ram_wvalid_272 && 0) begin
            write_burst_packed_done_277 <= 1;
          end 
          if(write_burst_block_ram_wvalid_272 && (write_burst_packed_length_276 <= 1)) begin
            write_burst_packed_fsm_49 <= write_burst_packed_fsm_49_init;
          end 
          if(write_burst_block_ram_wvalid_272 && 0) begin
            write_burst_packed_fsm_49 <= write_burst_packed_fsm_49_init;
          end 
          if(write_burst_block_ram_wquit_273) begin
            write_burst_packed_fsm_49 <= write_burst_packed_fsm_49_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_block_fsm_50_1 = 1;
  localparam write_burst_block_fsm_50_2 = 2;
  localparam write_burst_block_fsm_50_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_block_fsm_50 <= write_burst_block_fsm_50_init;
      write_burst_block_length_282 <= 0;
      write_burst_block_blocksize_283 <= 0;
      write_burst_block_done_284 <= 0;
      write_burst_block_count_285 <= 0;
    end else begin
      case(write_burst_block_fsm_50)
        write_burst_block_fsm_50_init: begin
          write_burst_block_length_282 <= _maxi_read_local_size_buf;
          write_burst_block_blocksize_283 <= _maxi_read_local_blocksize_buf;
          write_burst_block_done_284 <= 0;
          write_burst_block_count_285 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 5) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_block_fsm_50 <= write_burst_block_fsm_50_1;
          end 
        end
        write_burst_block_fsm_50_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_282 <= write_burst_block_length_282 - 1;
            write_burst_block_done_284 <= 0;
            write_burst_block_count_285 <= write_burst_block_count_285 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_282 <= 1)) begin
            write_burst_block_done_284 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_284 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_285 == write_burst_block_blocksize_283 - 1)) begin
            write_burst_block_count_285 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_285 == write_burst_block_blocksize_283 - 1)) begin
            write_burst_block_fsm_50 <= write_burst_block_fsm_50_2;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_282 <= 1)) begin
            write_burst_block_fsm_50 <= write_burst_block_fsm_50_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_50 <= write_burst_block_fsm_50_init;
          end 
          if(0) begin
            write_burst_block_fsm_50 <= write_burst_block_fsm_50_init;
          end 
        end
        write_burst_block_fsm_50_2: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_282 <= write_burst_block_length_282 - 1;
            write_burst_block_done_284 <= 0;
            write_burst_block_count_285 <= write_burst_block_count_285 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_282 <= 1)) begin
            write_burst_block_done_284 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_284 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_285 == write_burst_block_blocksize_283 - 1)) begin
            write_burst_block_count_285 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_285 == write_burst_block_blocksize_283 - 1)) begin
            write_burst_block_fsm_50 <= write_burst_block_fsm_50_3;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_282 <= 1)) begin
            write_burst_block_fsm_50 <= write_burst_block_fsm_50_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_50 <= write_burst_block_fsm_50_init;
          end 
          if(0) begin
            write_burst_block_fsm_50 <= write_burst_block_fsm_50_init;
          end 
        end
        write_burst_block_fsm_50_3: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_282 <= write_burst_block_length_282 - 1;
            write_burst_block_done_284 <= 0;
            write_burst_block_count_285 <= write_burst_block_count_285 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_282 <= 1)) begin
            write_burst_block_done_284 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_284 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_285 == write_burst_block_blocksize_283 - 1)) begin
            write_burst_block_count_285 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_285 == write_burst_block_blocksize_283 - 1)) begin
            write_burst_block_fsm_50 <= write_burst_block_fsm_50_1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_282 <= 1)) begin
            write_burst_block_fsm_50 <= write_burst_block_fsm_50_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_50 <= write_burst_block_fsm_50_init;
          end 
          if(0) begin
            write_burst_block_fsm_50 <= write_burst_block_fsm_50_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_51_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_51 <= write_burst_packed_fsm_51_init;
      write_burst_packed_addr_296 <= 0;
      write_burst_packed_stride_297 <= 0;
      write_burst_packed_length_298 <= 0;
      write_burst_packed_done_299 <= 0;
    end else begin
      case(write_burst_packed_fsm_51)
        write_burst_packed_fsm_51_init: begin
          write_burst_packed_addr_296 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_297 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_298 <= _maxi_read_local_size_buf;
          write_burst_packed_done_299 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 6) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_51 <= write_burst_packed_fsm_51_1;
          end 
        end
        write_burst_packed_fsm_51_1: begin
          if(write_burst_block_ram_wvalid_294) begin
            write_burst_packed_addr_296 <= write_burst_packed_addr_296 + write_burst_packed_stride_297;
            write_burst_packed_length_298 <= write_burst_packed_length_298 - 1;
            write_burst_packed_done_299 <= 0;
          end 
          if(write_burst_block_ram_wvalid_294 && (write_burst_packed_length_298 <= 1)) begin
            write_burst_packed_done_299 <= 1;
          end 
          if(write_burst_block_ram_wvalid_294 && 0) begin
            write_burst_packed_done_299 <= 1;
          end 
          if(write_burst_block_ram_wvalid_294 && (write_burst_packed_length_298 <= 1)) begin
            write_burst_packed_fsm_51 <= write_burst_packed_fsm_51_init;
          end 
          if(write_burst_block_ram_wvalid_294 && 0) begin
            write_burst_packed_fsm_51 <= write_burst_packed_fsm_51_init;
          end 
          if(write_burst_block_ram_wquit_295) begin
            write_burst_packed_fsm_51 <= write_burst_packed_fsm_51_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_52_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_52 <= write_burst_packed_fsm_52_init;
      write_burst_packed_addr_306 <= 0;
      write_burst_packed_stride_307 <= 0;
      write_burst_packed_length_308 <= 0;
      write_burst_packed_done_309 <= 0;
    end else begin
      case(write_burst_packed_fsm_52)
        write_burst_packed_fsm_52_init: begin
          write_burst_packed_addr_306 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_307 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_308 <= _maxi_read_local_size_buf;
          write_burst_packed_done_309 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 6) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_52 <= write_burst_packed_fsm_52_1;
          end 
        end
        write_burst_packed_fsm_52_1: begin
          if(write_burst_block_ram_wvalid_304) begin
            write_burst_packed_addr_306 <= write_burst_packed_addr_306 + write_burst_packed_stride_307;
            write_burst_packed_length_308 <= write_burst_packed_length_308 - 1;
            write_burst_packed_done_309 <= 0;
          end 
          if(write_burst_block_ram_wvalid_304 && (write_burst_packed_length_308 <= 1)) begin
            write_burst_packed_done_309 <= 1;
          end 
          if(write_burst_block_ram_wvalid_304 && 0) begin
            write_burst_packed_done_309 <= 1;
          end 
          if(write_burst_block_ram_wvalid_304 && (write_burst_packed_length_308 <= 1)) begin
            write_burst_packed_fsm_52 <= write_burst_packed_fsm_52_init;
          end 
          if(write_burst_block_ram_wvalid_304 && 0) begin
            write_burst_packed_fsm_52 <= write_burst_packed_fsm_52_init;
          end 
          if(write_burst_block_ram_wquit_305) begin
            write_burst_packed_fsm_52 <= write_burst_packed_fsm_52_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_53_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_53 <= write_burst_packed_fsm_53_init;
      write_burst_packed_addr_316 <= 0;
      write_burst_packed_stride_317 <= 0;
      write_burst_packed_length_318 <= 0;
      write_burst_packed_done_319 <= 0;
    end else begin
      case(write_burst_packed_fsm_53)
        write_burst_packed_fsm_53_init: begin
          write_burst_packed_addr_316 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_317 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_318 <= _maxi_read_local_size_buf;
          write_burst_packed_done_319 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 6) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_53 <= write_burst_packed_fsm_53_1;
          end 
        end
        write_burst_packed_fsm_53_1: begin
          if(write_burst_block_ram_wvalid_314) begin
            write_burst_packed_addr_316 <= write_burst_packed_addr_316 + write_burst_packed_stride_317;
            write_burst_packed_length_318 <= write_burst_packed_length_318 - 1;
            write_burst_packed_done_319 <= 0;
          end 
          if(write_burst_block_ram_wvalid_314 && (write_burst_packed_length_318 <= 1)) begin
            write_burst_packed_done_319 <= 1;
          end 
          if(write_burst_block_ram_wvalid_314 && 0) begin
            write_burst_packed_done_319 <= 1;
          end 
          if(write_burst_block_ram_wvalid_314 && (write_burst_packed_length_318 <= 1)) begin
            write_burst_packed_fsm_53 <= write_burst_packed_fsm_53_init;
          end 
          if(write_burst_block_ram_wvalid_314 && 0) begin
            write_burst_packed_fsm_53 <= write_burst_packed_fsm_53_init;
          end 
          if(write_burst_block_ram_wquit_315) begin
            write_burst_packed_fsm_53 <= write_burst_packed_fsm_53_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_block_fsm_54_1 = 1;
  localparam write_burst_block_fsm_54_2 = 2;
  localparam write_burst_block_fsm_54_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_block_fsm_54 <= write_burst_block_fsm_54_init;
      write_burst_block_length_324 <= 0;
      write_burst_block_blocksize_325 <= 0;
      write_burst_block_done_326 <= 0;
      write_burst_block_count_327 <= 0;
    end else begin
      case(write_burst_block_fsm_54)
        write_burst_block_fsm_54_init: begin
          write_burst_block_length_324 <= _maxi_read_local_size_buf;
          write_burst_block_blocksize_325 <= _maxi_read_local_blocksize_buf;
          write_burst_block_done_326 <= 0;
          write_burst_block_count_327 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 6) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_block_fsm_54 <= write_burst_block_fsm_54_1;
          end 
        end
        write_burst_block_fsm_54_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_324 <= write_burst_block_length_324 - 1;
            write_burst_block_done_326 <= 0;
            write_burst_block_count_327 <= write_burst_block_count_327 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_324 <= 1)) begin
            write_burst_block_done_326 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_326 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_327 == write_burst_block_blocksize_325 - 1)) begin
            write_burst_block_count_327 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_327 == write_burst_block_blocksize_325 - 1)) begin
            write_burst_block_fsm_54 <= write_burst_block_fsm_54_2;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_324 <= 1)) begin
            write_burst_block_fsm_54 <= write_burst_block_fsm_54_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_54 <= write_burst_block_fsm_54_init;
          end 
          if(0) begin
            write_burst_block_fsm_54 <= write_burst_block_fsm_54_init;
          end 
        end
        write_burst_block_fsm_54_2: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_324 <= write_burst_block_length_324 - 1;
            write_burst_block_done_326 <= 0;
            write_burst_block_count_327 <= write_burst_block_count_327 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_324 <= 1)) begin
            write_burst_block_done_326 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_326 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_327 == write_burst_block_blocksize_325 - 1)) begin
            write_burst_block_count_327 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_327 == write_burst_block_blocksize_325 - 1)) begin
            write_burst_block_fsm_54 <= write_burst_block_fsm_54_3;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_324 <= 1)) begin
            write_burst_block_fsm_54 <= write_burst_block_fsm_54_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_54 <= write_burst_block_fsm_54_init;
          end 
          if(0) begin
            write_burst_block_fsm_54 <= write_burst_block_fsm_54_init;
          end 
        end
        write_burst_block_fsm_54_3: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_block_length_324 <= write_burst_block_length_324 - 1;
            write_burst_block_done_326 <= 0;
            write_burst_block_count_327 <= write_burst_block_count_327 + 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_324 <= 1)) begin
            write_burst_block_done_326 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_done_326 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_327 == write_burst_block_blocksize_325 - 1)) begin
            write_burst_block_count_327 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_count_327 == write_burst_block_blocksize_325 - 1)) begin
            write_burst_block_fsm_54 <= write_burst_block_fsm_54_1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_block_length_324 <= 1)) begin
            write_burst_block_fsm_54 <= write_burst_block_fsm_54_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_block_fsm_54 <= write_burst_block_fsm_54_init;
          end 
          if(0) begin
            write_burst_block_fsm_54 <= write_burst_block_fsm_54_init;
          end 
        end
      endcase
    end
  end

  localparam conv2d_4_comp_fsm_1 = 1;
  localparam conv2d_4_comp_fsm_2 = 2;
  localparam conv2d_4_comp_fsm_3 = 3;
  localparam conv2d_4_comp_fsm_4 = 4;
  localparam conv2d_4_comp_fsm_5 = 5;
  localparam conv2d_4_comp_fsm_6 = 6;

  always @(posedge CLK) begin
    if(RST) begin
      conv2d_4_comp_fsm <= conv2d_4_comp_fsm_init;
      conv2d_4_stream_act_local_0 <= 0;
      conv2d_4_stream_act_local_1 <= 0;
      conv2d_4_stream_act_local_2 <= 0;
      conv2d_4_stream_act_local_3 <= 0;
      conv2d_4_stream_act_local_4 <= 0;
      conv2d_4_stream_act_local_5 <= 0;
      conv2d_4_stream_act_local_6 <= 0;
      conv2d_4_stream_act_local_7 <= 0;
      conv2d_4_stream_act_local_8 <= 0;
      conv2d_4_stream_out_local_col <= 0;
      conv2d_4_stream_out_local_val <= 0;
      conv2d_4_col_count <= 0;
      conv2d_4_col_select <= 0;
      conv2d_4_filter_page_comp_offset_buf <= 0;
      conv2d_4_act_page_comp_offset_buf_0 <= 0;
      conv2d_4_act_page_comp_offset_buf_1 <= 0;
      conv2d_4_act_page_comp_offset_buf_2 <= 0;
      conv2d_4_out_page_comp_offset_buf <= 0;
      conv2d_4_row_count_buf <= 0;
      conv2d_4_row_select_buf <= 0;
      conv2d_4_och_count_buf <= 0;
      conv2d_4_next_stream_num_ops <= 0;
      conv2d_4_stream_pad_masks <= 0;
      conv2d_4_sync_comp_count <= 0;
    end else begin
      if(_stream_conv2d_4_sink_stop) begin
        conv2d_4_sync_comp_count <= conv2d_4_sync_comp_count + 1;
      end 
      if(control_conv2d_4 == 6) begin
        conv2d_4_sync_comp_count <= 0;
      end 
      case(conv2d_4_comp_fsm)
        conv2d_4_comp_fsm_init: begin
          if((control_conv2d_4 == 25) && !conv2d_4_skip_comp) begin
            conv2d_4_comp_fsm <= conv2d_4_comp_fsm_1;
          end 
        end
        conv2d_4_comp_fsm_1: begin
          conv2d_4_stream_act_local_0 <= 0;
          if(cparam_conv2d_4_stream_act_local_small_flags_0) begin
            conv2d_4_stream_act_local_0 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_4_stream_act_local_large_flags_0) begin
            conv2d_4_stream_act_local_0 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          conv2d_4_stream_act_local_1 <= 0;
          if(cparam_conv2d_4_stream_act_local_small_flags_1) begin
            conv2d_4_stream_act_local_1 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_4_stream_act_local_large_flags_1) begin
            conv2d_4_stream_act_local_1 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          conv2d_4_stream_act_local_2 <= 0;
          if(cparam_conv2d_4_stream_act_local_small_flags_2) begin
            conv2d_4_stream_act_local_2 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_4_stream_act_local_large_flags_2) begin
            conv2d_4_stream_act_local_2 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          conv2d_4_stream_act_local_3 <= 0;
          if(cparam_conv2d_4_stream_act_local_small_flags_0) begin
            conv2d_4_stream_act_local_3 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_4_stream_act_local_large_flags_0) begin
            conv2d_4_stream_act_local_3 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          conv2d_4_stream_act_local_4 <= 0;
          if(cparam_conv2d_4_stream_act_local_small_flags_1) begin
            conv2d_4_stream_act_local_4 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_4_stream_act_local_large_flags_1) begin
            conv2d_4_stream_act_local_4 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          conv2d_4_stream_act_local_5 <= 0;
          if(cparam_conv2d_4_stream_act_local_small_flags_2) begin
            conv2d_4_stream_act_local_5 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_4_stream_act_local_large_flags_2) begin
            conv2d_4_stream_act_local_5 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          conv2d_4_stream_act_local_6 <= 0;
          if(cparam_conv2d_4_stream_act_local_small_flags_0) begin
            conv2d_4_stream_act_local_6 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_4_stream_act_local_large_flags_0) begin
            conv2d_4_stream_act_local_6 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          conv2d_4_stream_act_local_7 <= 0;
          if(cparam_conv2d_4_stream_act_local_small_flags_1) begin
            conv2d_4_stream_act_local_7 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_4_stream_act_local_large_flags_1) begin
            conv2d_4_stream_act_local_7 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          conv2d_4_stream_act_local_8 <= 0;
          if(cparam_conv2d_4_stream_act_local_small_flags_2) begin
            conv2d_4_stream_act_local_8 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if(cparam_conv2d_4_stream_act_local_large_flags_2) begin
            conv2d_4_stream_act_local_8 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          conv2d_4_stream_out_local_col <= 0;
          if((cparam_conv2d_4_data_stationary == 1) && (conv2d_4_och_count == 0)) begin
            conv2d_4_stream_out_local_val <= 0;
          end 
          conv2d_4_col_count <= 0;
          conv2d_4_col_select <= cparam_conv2d_4_col_select_initval;
          conv2d_4_filter_page_comp_offset_buf <= conv2d_4_filter_page_comp_offset;
          conv2d_4_act_page_comp_offset_buf_0 <= conv2d_4_act_page_comp_offset_0;
          conv2d_4_act_page_comp_offset_buf_1 <= conv2d_4_act_page_comp_offset_1;
          conv2d_4_act_page_comp_offset_buf_2 <= conv2d_4_act_page_comp_offset_2;
          conv2d_4_out_page_comp_offset_buf <= conv2d_4_out_page_comp_offset;
          conv2d_4_row_count_buf <= conv2d_4_row_count;
          conv2d_4_row_select_buf <= conv2d_4_row_select;
          conv2d_4_och_count_buf <= conv2d_4_och_count;
          conv2d_4_next_stream_num_ops <= (conv2d_4_och_count >= cparam_conv2d_4_max_och_count)? cparam_conv2d_4_stream_num_ops_res : cparam_conv2d_4_stream_num_ops;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_2;
        end
        conv2d_4_comp_fsm_2: begin
          conv2d_4_stream_pad_masks <= { conv2d_4_stream_pad_mask_2_2, conv2d_4_stream_pad_mask_2_1, conv2d_4_stream_pad_mask_2_0, conv2d_4_stream_pad_mask_1_2, conv2d_4_stream_pad_mask_1_1, conv2d_4_stream_pad_mask_1_0, conv2d_4_stream_pad_mask_0_2, conv2d_4_stream_pad_mask_0_1, conv2d_4_stream_pad_mask_0_0 };
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_3;
        end
        conv2d_4_comp_fsm_3: begin
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          if(_stream_conv2d_4_stream_oready) begin
            conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
          end 
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_4;
        end
        conv2d_4_comp_fsm_4: begin
          if(!_stream_conv2d_4_source_busy) begin
            conv2d_4_comp_fsm <= conv2d_4_comp_fsm_5;
          end 
        end
        conv2d_4_comp_fsm_5: begin
          if(_stream_conv2d_4_busy) begin
            conv2d_4_comp_fsm <= conv2d_4_comp_fsm_6;
          end 
        end
        conv2d_4_comp_fsm_6: begin
          if(!((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_0 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_1 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_2 : 0)) begin
            conv2d_4_stream_act_local_0 <= conv2d_4_stream_act_local_0 + cparam_conv2d_4_inc_act_laddr_small;
          end 
          if((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_0 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_1 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_2 : 0) begin
            conv2d_4_stream_act_local_0 <= conv2d_4_stream_act_local_0 + cparam_conv2d_4_inc_act_laddr_large;
          end 
          if(conv2d_4_col_count >= cparam_conv2d_4_max_col_count) begin
            conv2d_4_stream_act_local_0 <= 0;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_small_flags_0) begin
            conv2d_4_stream_act_local_0 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_large_flags_0) begin
            conv2d_4_stream_act_local_0 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          if(!((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_3 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_4 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_5 : 0)) begin
            conv2d_4_stream_act_local_1 <= conv2d_4_stream_act_local_1 + cparam_conv2d_4_inc_act_laddr_small;
          end 
          if((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_3 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_4 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_5 : 0) begin
            conv2d_4_stream_act_local_1 <= conv2d_4_stream_act_local_1 + cparam_conv2d_4_inc_act_laddr_large;
          end 
          if(conv2d_4_col_count >= cparam_conv2d_4_max_col_count) begin
            conv2d_4_stream_act_local_1 <= 0;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_small_flags_1) begin
            conv2d_4_stream_act_local_1 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_large_flags_1) begin
            conv2d_4_stream_act_local_1 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          if(!((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_6 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_7 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_8 : 0)) begin
            conv2d_4_stream_act_local_2 <= conv2d_4_stream_act_local_2 + cparam_conv2d_4_inc_act_laddr_small;
          end 
          if((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_6 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_7 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_8 : 0) begin
            conv2d_4_stream_act_local_2 <= conv2d_4_stream_act_local_2 + cparam_conv2d_4_inc_act_laddr_large;
          end 
          if(conv2d_4_col_count >= cparam_conv2d_4_max_col_count) begin
            conv2d_4_stream_act_local_2 <= 0;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_small_flags_2) begin
            conv2d_4_stream_act_local_2 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_large_flags_2) begin
            conv2d_4_stream_act_local_2 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          if(!((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_9 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_10 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_11 : 0)) begin
            conv2d_4_stream_act_local_3 <= conv2d_4_stream_act_local_3 + cparam_conv2d_4_inc_act_laddr_small;
          end 
          if((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_9 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_10 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_11 : 0) begin
            conv2d_4_stream_act_local_3 <= conv2d_4_stream_act_local_3 + cparam_conv2d_4_inc_act_laddr_large;
          end 
          if(conv2d_4_col_count >= cparam_conv2d_4_max_col_count) begin
            conv2d_4_stream_act_local_3 <= 0;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_small_flags_0) begin
            conv2d_4_stream_act_local_3 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_large_flags_0) begin
            conv2d_4_stream_act_local_3 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          if(!((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_12 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_13 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_14 : 0)) begin
            conv2d_4_stream_act_local_4 <= conv2d_4_stream_act_local_4 + cparam_conv2d_4_inc_act_laddr_small;
          end 
          if((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_12 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_13 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_14 : 0) begin
            conv2d_4_stream_act_local_4 <= conv2d_4_stream_act_local_4 + cparam_conv2d_4_inc_act_laddr_large;
          end 
          if(conv2d_4_col_count >= cparam_conv2d_4_max_col_count) begin
            conv2d_4_stream_act_local_4 <= 0;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_small_flags_1) begin
            conv2d_4_stream_act_local_4 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_large_flags_1) begin
            conv2d_4_stream_act_local_4 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          if(!((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_15 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_16 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_17 : 0)) begin
            conv2d_4_stream_act_local_5 <= conv2d_4_stream_act_local_5 + cparam_conv2d_4_inc_act_laddr_small;
          end 
          if((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_15 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_16 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_17 : 0) begin
            conv2d_4_stream_act_local_5 <= conv2d_4_stream_act_local_5 + cparam_conv2d_4_inc_act_laddr_large;
          end 
          if(conv2d_4_col_count >= cparam_conv2d_4_max_col_count) begin
            conv2d_4_stream_act_local_5 <= 0;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_small_flags_2) begin
            conv2d_4_stream_act_local_5 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_large_flags_2) begin
            conv2d_4_stream_act_local_5 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          if(!((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_18 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_19 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_20 : 0)) begin
            conv2d_4_stream_act_local_6 <= conv2d_4_stream_act_local_6 + cparam_conv2d_4_inc_act_laddr_small;
          end 
          if((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_18 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_19 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_20 : 0) begin
            conv2d_4_stream_act_local_6 <= conv2d_4_stream_act_local_6 + cparam_conv2d_4_inc_act_laddr_large;
          end 
          if(conv2d_4_col_count >= cparam_conv2d_4_max_col_count) begin
            conv2d_4_stream_act_local_6 <= 0;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_small_flags_0) begin
            conv2d_4_stream_act_local_6 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_large_flags_0) begin
            conv2d_4_stream_act_local_6 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          if(!((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_21 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_22 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_23 : 0)) begin
            conv2d_4_stream_act_local_7 <= conv2d_4_stream_act_local_7 + cparam_conv2d_4_inc_act_laddr_small;
          end 
          if((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_21 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_22 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_23 : 0) begin
            conv2d_4_stream_act_local_7 <= conv2d_4_stream_act_local_7 + cparam_conv2d_4_inc_act_laddr_large;
          end 
          if(conv2d_4_col_count >= cparam_conv2d_4_max_col_count) begin
            conv2d_4_stream_act_local_7 <= 0;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_small_flags_1) begin
            conv2d_4_stream_act_local_7 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_large_flags_1) begin
            conv2d_4_stream_act_local_7 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          if(!((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_24 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_25 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_26 : 0)) begin
            conv2d_4_stream_act_local_8 <= conv2d_4_stream_act_local_8 + cparam_conv2d_4_inc_act_laddr_small;
          end 
          if((conv2d_4_col_select == 0)? cparam_conv2d_4_inc_act_laddr_conds_24 : 
          (conv2d_4_col_select == 1)? cparam_conv2d_4_inc_act_laddr_conds_25 : 
          (conv2d_4_col_select == 2)? cparam_conv2d_4_inc_act_laddr_conds_26 : 0) begin
            conv2d_4_stream_act_local_8 <= conv2d_4_stream_act_local_8 + cparam_conv2d_4_inc_act_laddr_large;
          end 
          if(conv2d_4_col_count >= cparam_conv2d_4_max_col_count) begin
            conv2d_4_stream_act_local_8 <= 0;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_small_flags_2) begin
            conv2d_4_stream_act_local_8 <= cparam_conv2d_4_stream_act_local_small_offset;
          end 
          if((conv2d_4_col_count >= cparam_conv2d_4_max_col_count) && cparam_conv2d_4_stream_act_local_large_flags_2) begin
            conv2d_4_stream_act_local_8 <= cparam_conv2d_4_stream_act_local_large_offset;
          end 
          if(cparam_conv2d_4_data_stationary == 0) begin
            conv2d_4_stream_out_local_col <= conv2d_4_stream_out_local_col + conv2d_4_next_stream_num_ops;
          end 
          if((cparam_conv2d_4_data_stationary == 0) && (conv2d_4_col_count >= cparam_conv2d_4_max_col_count)) begin
            conv2d_4_stream_out_local_col <= 0;
          end 
          if(cparam_conv2d_4_data_stationary == 1) begin
            conv2d_4_stream_out_local_col <= conv2d_4_stream_out_local_col + cparam_conv2d_4_inc_out_laddr_col;
          end 
          if((cparam_conv2d_4_data_stationary == 1) && (conv2d_4_col_count >= cparam_conv2d_4_max_col_count)) begin
            conv2d_4_stream_out_local_val <= conv2d_4_stream_out_local_val + conv2d_4_next_stream_num_ops;
            conv2d_4_stream_out_local_col <= 0;
          end 
          conv2d_4_col_count <= conv2d_4_col_count + cparam_conv2d_4_stride_col_par_col;
          if(conv2d_4_col_count >= cparam_conv2d_4_max_col_count) begin
            conv2d_4_col_count <= 0;
          end 
          conv2d_4_col_select <= conv2d_4_col_select + cparam_conv2d_4_stride_col_mod_filter_num;
          if(conv2d_4_col_select + cparam_conv2d_4_stride_col_mod_filter_num >= 3) begin
            conv2d_4_col_select <= conv2d_4_col_select - cparam_conv2d_4_filter_num_col_minus_stride_col_mod;
          end 
          if(conv2d_4_col_count >= cparam_conv2d_4_max_col_count) begin
            conv2d_4_col_select <= cparam_conv2d_4_col_select_initval;
          end 
          conv2d_4_comp_fsm <= conv2d_4_comp_fsm_2;
          if(conv2d_4_col_count >= cparam_conv2d_4_max_col_count) begin
            conv2d_4_comp_fsm <= conv2d_4_comp_fsm_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_336 <= 0;
    end else begin
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_7_source_ram_renable && (_stream_conv2d_4_source_7_source_sel == 1)) begin
        _tmp_336 <= read_rtl_bank_335;
      end 
    end
  end

  localparam _stream_conv2d_4_source_7_source_pat_fsm_0_1 = 1;
  localparam _stream_conv2d_4_source_7_source_pat_fsm_0_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_7_source_pat_fsm_0 <= _stream_conv2d_4_source_7_source_pat_fsm_0_init;
    end else begin
      case(_stream_conv2d_4_source_7_source_pat_fsm_0)
        _stream_conv2d_4_source_7_source_pat_fsm_0_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_7_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_7_source_pat_fsm_0 <= _stream_conv2d_4_source_7_source_pat_fsm_0_1;
          end 
        end
        _stream_conv2d_4_source_7_source_pat_fsm_0_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_7_source_pat_fsm_0 <= _stream_conv2d_4_source_7_source_pat_fsm_0_init;
          end 
          if((_source_stream_conv2d_4_source_7_pat_count_0 == 0) && (_source_stream_conv2d_4_source_7_pat_count_1 == 0) && (_source_stream_conv2d_4_source_7_pat_count_2 == 0) && (_source_stream_conv2d_4_source_7_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_7_source_pat_fsm_0 <= _stream_conv2d_4_source_7_source_pat_fsm_0_2;
          end 
        end
        _stream_conv2d_4_source_7_source_pat_fsm_0_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_7_source_pat_fsm_0 <= _stream_conv2d_4_source_7_source_pat_fsm_0_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_346 <= 0;
    end else begin
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_9_source_ram_renable && (_stream_conv2d_4_source_9_source_sel == 2)) begin
        _tmp_346 <= read_rtl_bank_345;
      end 
    end
  end

  localparam _stream_conv2d_4_source_9_source_pat_fsm_1_1 = 1;
  localparam _stream_conv2d_4_source_9_source_pat_fsm_1_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_9_source_pat_fsm_1 <= _stream_conv2d_4_source_9_source_pat_fsm_1_init;
    end else begin
      case(_stream_conv2d_4_source_9_source_pat_fsm_1)
        _stream_conv2d_4_source_9_source_pat_fsm_1_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_9_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_9_source_pat_fsm_1 <= _stream_conv2d_4_source_9_source_pat_fsm_1_1;
          end 
        end
        _stream_conv2d_4_source_9_source_pat_fsm_1_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_9_source_pat_fsm_1 <= _stream_conv2d_4_source_9_source_pat_fsm_1_init;
          end 
          if((_source_stream_conv2d_4_source_9_pat_count_0 == 0) && (_source_stream_conv2d_4_source_9_pat_count_1 == 0) && (_source_stream_conv2d_4_source_9_pat_count_2 == 0) && (_source_stream_conv2d_4_source_9_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_9_source_pat_fsm_1 <= _stream_conv2d_4_source_9_source_pat_fsm_1_2;
          end 
        end
        _stream_conv2d_4_source_9_source_pat_fsm_1_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_9_source_pat_fsm_1 <= _stream_conv2d_4_source_9_source_pat_fsm_1_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_365 <= 0;
    end else begin
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_20_source_ram_renable && (_stream_conv2d_4_source_20_source_sel == 3)) begin
        _tmp_365 <= read_rtl_bank_364;
      end 
    end
  end

  localparam _stream_conv2d_4_source_20_source_pat_fsm_2_1 = 1;
  localparam _stream_conv2d_4_source_20_source_pat_fsm_2_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_20_source_pat_fsm_2 <= _stream_conv2d_4_source_20_source_pat_fsm_2_init;
    end else begin
      case(_stream_conv2d_4_source_20_source_pat_fsm_2)
        _stream_conv2d_4_source_20_source_pat_fsm_2_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_20_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_20_source_pat_fsm_2 <= _stream_conv2d_4_source_20_source_pat_fsm_2_1;
          end 
        end
        _stream_conv2d_4_source_20_source_pat_fsm_2_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_20_source_pat_fsm_2 <= _stream_conv2d_4_source_20_source_pat_fsm_2_init;
          end 
          if((_source_stream_conv2d_4_source_20_pat_count_0 == 0) && (_source_stream_conv2d_4_source_20_pat_count_1 == 0) && (_source_stream_conv2d_4_source_20_pat_count_2 == 0) && (_source_stream_conv2d_4_source_20_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_20_source_pat_fsm_2 <= _stream_conv2d_4_source_20_source_pat_fsm_2_2;
          end 
        end
        _stream_conv2d_4_source_20_source_pat_fsm_2_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_20_source_pat_fsm_2 <= _stream_conv2d_4_source_20_source_pat_fsm_2_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_374 <= 0;
    end else begin
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_21_source_ram_renable && (_stream_conv2d_4_source_21_source_sel == 4)) begin
        _tmp_374 <= read_rtl_bank_373;
      end 
    end
  end

  localparam _stream_conv2d_4_source_21_source_pat_fsm_3_1 = 1;
  localparam _stream_conv2d_4_source_21_source_pat_fsm_3_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_21_source_pat_fsm_3 <= _stream_conv2d_4_source_21_source_pat_fsm_3_init;
    end else begin
      case(_stream_conv2d_4_source_21_source_pat_fsm_3)
        _stream_conv2d_4_source_21_source_pat_fsm_3_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_21_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_21_source_pat_fsm_3 <= _stream_conv2d_4_source_21_source_pat_fsm_3_1;
          end 
        end
        _stream_conv2d_4_source_21_source_pat_fsm_3_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_21_source_pat_fsm_3 <= _stream_conv2d_4_source_21_source_pat_fsm_3_init;
          end 
          if((_source_stream_conv2d_4_source_21_pat_count_0 == 0) && (_source_stream_conv2d_4_source_21_pat_count_1 == 0) && (_source_stream_conv2d_4_source_21_pat_count_2 == 0) && (_source_stream_conv2d_4_source_21_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_21_source_pat_fsm_3 <= _stream_conv2d_4_source_21_source_pat_fsm_3_2;
          end 
        end
        _stream_conv2d_4_source_21_source_pat_fsm_3_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_21_source_pat_fsm_3 <= _stream_conv2d_4_source_21_source_pat_fsm_3_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_383 <= 0;
    end else begin
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_22_source_ram_renable && (_stream_conv2d_4_source_22_source_sel == 5)) begin
        _tmp_383 <= read_rtl_bank_382;
      end 
    end
  end

  localparam _stream_conv2d_4_source_22_source_pat_fsm_4_1 = 1;
  localparam _stream_conv2d_4_source_22_source_pat_fsm_4_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_22_source_pat_fsm_4 <= _stream_conv2d_4_source_22_source_pat_fsm_4_init;
    end else begin
      case(_stream_conv2d_4_source_22_source_pat_fsm_4)
        _stream_conv2d_4_source_22_source_pat_fsm_4_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_22_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_22_source_pat_fsm_4 <= _stream_conv2d_4_source_22_source_pat_fsm_4_1;
          end 
        end
        _stream_conv2d_4_source_22_source_pat_fsm_4_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_22_source_pat_fsm_4 <= _stream_conv2d_4_source_22_source_pat_fsm_4_init;
          end 
          if((_source_stream_conv2d_4_source_22_pat_count_0 == 0) && (_source_stream_conv2d_4_source_22_pat_count_1 == 0) && (_source_stream_conv2d_4_source_22_pat_count_2 == 0) && (_source_stream_conv2d_4_source_22_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_22_source_pat_fsm_4 <= _stream_conv2d_4_source_22_source_pat_fsm_4_2;
          end 
        end
        _stream_conv2d_4_source_22_source_pat_fsm_4_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_22_source_pat_fsm_4 <= _stream_conv2d_4_source_22_source_pat_fsm_4_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_392 <= 0;
    end else begin
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_23_source_ram_renable && (_stream_conv2d_4_source_23_source_sel == 6)) begin
        _tmp_392 <= read_rtl_bank_391;
      end 
    end
  end

  localparam _stream_conv2d_4_source_23_source_pat_fsm_5_1 = 1;
  localparam _stream_conv2d_4_source_23_source_pat_fsm_5_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_23_source_pat_fsm_5 <= _stream_conv2d_4_source_23_source_pat_fsm_5_init;
    end else begin
      case(_stream_conv2d_4_source_23_source_pat_fsm_5)
        _stream_conv2d_4_source_23_source_pat_fsm_5_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_23_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_23_source_pat_fsm_5 <= _stream_conv2d_4_source_23_source_pat_fsm_5_1;
          end 
        end
        _stream_conv2d_4_source_23_source_pat_fsm_5_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_23_source_pat_fsm_5 <= _stream_conv2d_4_source_23_source_pat_fsm_5_init;
          end 
          if((_source_stream_conv2d_4_source_23_pat_count_0 == 0) && (_source_stream_conv2d_4_source_23_pat_count_1 == 0) && (_source_stream_conv2d_4_source_23_pat_count_2 == 0) && (_source_stream_conv2d_4_source_23_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_23_source_pat_fsm_5 <= _stream_conv2d_4_source_23_source_pat_fsm_5_2;
          end 
        end
        _stream_conv2d_4_source_23_source_pat_fsm_5_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_23_source_pat_fsm_5 <= _stream_conv2d_4_source_23_source_pat_fsm_5_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_401 <= 0;
    end else begin
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_24_source_ram_renable && (_stream_conv2d_4_source_24_source_sel == 7)) begin
        _tmp_401 <= read_rtl_bank_400;
      end 
    end
  end

  localparam _stream_conv2d_4_source_24_source_pat_fsm_6_1 = 1;
  localparam _stream_conv2d_4_source_24_source_pat_fsm_6_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_24_source_pat_fsm_6 <= _stream_conv2d_4_source_24_source_pat_fsm_6_init;
    end else begin
      case(_stream_conv2d_4_source_24_source_pat_fsm_6)
        _stream_conv2d_4_source_24_source_pat_fsm_6_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_24_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_24_source_pat_fsm_6 <= _stream_conv2d_4_source_24_source_pat_fsm_6_1;
          end 
        end
        _stream_conv2d_4_source_24_source_pat_fsm_6_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_24_source_pat_fsm_6 <= _stream_conv2d_4_source_24_source_pat_fsm_6_init;
          end 
          if((_source_stream_conv2d_4_source_24_pat_count_0 == 0) && (_source_stream_conv2d_4_source_24_pat_count_1 == 0) && (_source_stream_conv2d_4_source_24_pat_count_2 == 0) && (_source_stream_conv2d_4_source_24_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_24_source_pat_fsm_6 <= _stream_conv2d_4_source_24_source_pat_fsm_6_2;
          end 
        end
        _stream_conv2d_4_source_24_source_pat_fsm_6_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_24_source_pat_fsm_6 <= _stream_conv2d_4_source_24_source_pat_fsm_6_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_410 <= 0;
    end else begin
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_25_source_ram_renable && (_stream_conv2d_4_source_25_source_sel == 8)) begin
        _tmp_410 <= read_rtl_bank_409;
      end 
    end
  end

  localparam _stream_conv2d_4_source_25_source_pat_fsm_7_1 = 1;
  localparam _stream_conv2d_4_source_25_source_pat_fsm_7_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_25_source_pat_fsm_7 <= _stream_conv2d_4_source_25_source_pat_fsm_7_init;
    end else begin
      case(_stream_conv2d_4_source_25_source_pat_fsm_7)
        _stream_conv2d_4_source_25_source_pat_fsm_7_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_25_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_25_source_pat_fsm_7 <= _stream_conv2d_4_source_25_source_pat_fsm_7_1;
          end 
        end
        _stream_conv2d_4_source_25_source_pat_fsm_7_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_25_source_pat_fsm_7 <= _stream_conv2d_4_source_25_source_pat_fsm_7_init;
          end 
          if((_source_stream_conv2d_4_source_25_pat_count_0 == 0) && (_source_stream_conv2d_4_source_25_pat_count_1 == 0) && (_source_stream_conv2d_4_source_25_pat_count_2 == 0) && (_source_stream_conv2d_4_source_25_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_25_source_pat_fsm_7 <= _stream_conv2d_4_source_25_source_pat_fsm_7_2;
          end 
        end
        _stream_conv2d_4_source_25_source_pat_fsm_7_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_25_source_pat_fsm_7 <= _stream_conv2d_4_source_25_source_pat_fsm_7_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_419 <= 0;
    end else begin
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_26_source_ram_renable && (_stream_conv2d_4_source_26_source_sel == 9)) begin
        _tmp_419 <= read_rtl_bank_418;
      end 
    end
  end

  localparam _stream_conv2d_4_source_26_source_pat_fsm_8_1 = 1;
  localparam _stream_conv2d_4_source_26_source_pat_fsm_8_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_26_source_pat_fsm_8 <= _stream_conv2d_4_source_26_source_pat_fsm_8_init;
    end else begin
      case(_stream_conv2d_4_source_26_source_pat_fsm_8)
        _stream_conv2d_4_source_26_source_pat_fsm_8_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_26_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_26_source_pat_fsm_8 <= _stream_conv2d_4_source_26_source_pat_fsm_8_1;
          end 
        end
        _stream_conv2d_4_source_26_source_pat_fsm_8_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_26_source_pat_fsm_8 <= _stream_conv2d_4_source_26_source_pat_fsm_8_init;
          end 
          if((_source_stream_conv2d_4_source_26_pat_count_0 == 0) && (_source_stream_conv2d_4_source_26_pat_count_1 == 0) && (_source_stream_conv2d_4_source_26_pat_count_2 == 0) && (_source_stream_conv2d_4_source_26_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_26_source_pat_fsm_8 <= _stream_conv2d_4_source_26_source_pat_fsm_8_2;
          end 
        end
        _stream_conv2d_4_source_26_source_pat_fsm_8_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_26_source_pat_fsm_8 <= _stream_conv2d_4_source_26_source_pat_fsm_8_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_428 <= 0;
    end else begin
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_27_source_ram_renable && (_stream_conv2d_4_source_27_source_sel == 10)) begin
        _tmp_428 <= read_rtl_bank_427;
      end 
    end
  end

  localparam _stream_conv2d_4_source_27_source_pat_fsm_9_1 = 1;
  localparam _stream_conv2d_4_source_27_source_pat_fsm_9_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_27_source_pat_fsm_9 <= _stream_conv2d_4_source_27_source_pat_fsm_9_init;
    end else begin
      case(_stream_conv2d_4_source_27_source_pat_fsm_9)
        _stream_conv2d_4_source_27_source_pat_fsm_9_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_27_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_27_source_pat_fsm_9 <= _stream_conv2d_4_source_27_source_pat_fsm_9_1;
          end 
        end
        _stream_conv2d_4_source_27_source_pat_fsm_9_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_27_source_pat_fsm_9 <= _stream_conv2d_4_source_27_source_pat_fsm_9_init;
          end 
          if((_source_stream_conv2d_4_source_27_pat_count_0 == 0) && (_source_stream_conv2d_4_source_27_pat_count_1 == 0) && (_source_stream_conv2d_4_source_27_pat_count_2 == 0) && (_source_stream_conv2d_4_source_27_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_27_source_pat_fsm_9 <= _stream_conv2d_4_source_27_source_pat_fsm_9_2;
          end 
        end
        _stream_conv2d_4_source_27_source_pat_fsm_9_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_27_source_pat_fsm_9 <= _stream_conv2d_4_source_27_source_pat_fsm_9_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_437 <= 0;
    end else begin
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_28_source_ram_renable && (_stream_conv2d_4_source_28_source_sel == 11)) begin
        _tmp_437 <= read_rtl_bank_436;
      end 
    end
  end

  localparam _stream_conv2d_4_source_28_source_pat_fsm_10_1 = 1;
  localparam _stream_conv2d_4_source_28_source_pat_fsm_10_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_28_source_pat_fsm_10 <= _stream_conv2d_4_source_28_source_pat_fsm_10_init;
    end else begin
      case(_stream_conv2d_4_source_28_source_pat_fsm_10)
        _stream_conv2d_4_source_28_source_pat_fsm_10_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_28_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_28_source_pat_fsm_10 <= _stream_conv2d_4_source_28_source_pat_fsm_10_1;
          end 
        end
        _stream_conv2d_4_source_28_source_pat_fsm_10_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_28_source_pat_fsm_10 <= _stream_conv2d_4_source_28_source_pat_fsm_10_init;
          end 
          if((_source_stream_conv2d_4_source_28_pat_count_0 == 0) && (_source_stream_conv2d_4_source_28_pat_count_1 == 0) && (_source_stream_conv2d_4_source_28_pat_count_2 == 0) && (_source_stream_conv2d_4_source_28_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_28_source_pat_fsm_10 <= _stream_conv2d_4_source_28_source_pat_fsm_10_2;
          end 
        end
        _stream_conv2d_4_source_28_source_pat_fsm_10_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_28_source_pat_fsm_10 <= _stream_conv2d_4_source_28_source_pat_fsm_10_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_446 <= 0;
    end else begin
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_29_source_ram_renable && (_stream_conv2d_4_source_29_source_sel == 12)) begin
        _tmp_446 <= read_rtl_bank_445;
      end 
    end
  end

  localparam _stream_conv2d_4_source_29_source_pat_fsm_11_1 = 1;
  localparam _stream_conv2d_4_source_29_source_pat_fsm_11_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_29_source_pat_fsm_11 <= _stream_conv2d_4_source_29_source_pat_fsm_11_init;
    end else begin
      case(_stream_conv2d_4_source_29_source_pat_fsm_11)
        _stream_conv2d_4_source_29_source_pat_fsm_11_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_29_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_29_source_pat_fsm_11 <= _stream_conv2d_4_source_29_source_pat_fsm_11_1;
          end 
        end
        _stream_conv2d_4_source_29_source_pat_fsm_11_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_29_source_pat_fsm_11 <= _stream_conv2d_4_source_29_source_pat_fsm_11_init;
          end 
          if((_source_stream_conv2d_4_source_29_pat_count_0 == 0) && (_source_stream_conv2d_4_source_29_pat_count_1 == 0) && (_source_stream_conv2d_4_source_29_pat_count_2 == 0) && (_source_stream_conv2d_4_source_29_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_29_source_pat_fsm_11 <= _stream_conv2d_4_source_29_source_pat_fsm_11_2;
          end 
        end
        _stream_conv2d_4_source_29_source_pat_fsm_11_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_29_source_pat_fsm_11 <= _stream_conv2d_4_source_29_source_pat_fsm_11_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_455 <= 0;
      _tmp_1364 <= 0;
    end else begin
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_30_source_ram_renable && (_stream_conv2d_4_source_30_source_sel == 13)) begin
        _tmp_455 <= read_rtl_bank_454;
      end 
      if(_stream_matmul_11_stream_oready && _stream_matmul_11_source_7_source_ram_renable && (_stream_matmul_11_source_7_source_sel == 1)) begin
        _tmp_1364 <= read_rtl_bank_1363;
      end 
    end
  end

  localparam _stream_conv2d_4_source_30_source_pat_fsm_12_1 = 1;
  localparam _stream_conv2d_4_source_30_source_pat_fsm_12_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_30_source_pat_fsm_12 <= _stream_conv2d_4_source_30_source_pat_fsm_12_init;
    end else begin
      case(_stream_conv2d_4_source_30_source_pat_fsm_12)
        _stream_conv2d_4_source_30_source_pat_fsm_12_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_30_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_30_source_pat_fsm_12 <= _stream_conv2d_4_source_30_source_pat_fsm_12_1;
          end 
        end
        _stream_conv2d_4_source_30_source_pat_fsm_12_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_30_source_pat_fsm_12 <= _stream_conv2d_4_source_30_source_pat_fsm_12_init;
          end 
          if((_source_stream_conv2d_4_source_30_pat_count_0 == 0) && (_source_stream_conv2d_4_source_30_pat_count_1 == 0) && (_source_stream_conv2d_4_source_30_pat_count_2 == 0) && (_source_stream_conv2d_4_source_30_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_30_source_pat_fsm_12 <= _stream_conv2d_4_source_30_source_pat_fsm_12_2;
          end 
        end
        _stream_conv2d_4_source_30_source_pat_fsm_12_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_30_source_pat_fsm_12 <= _stream_conv2d_4_source_30_source_pat_fsm_12_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_464 <= 0;
      _tmp_1374 <= 0;
    end else begin
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_31_source_ram_renable && (_stream_conv2d_4_source_31_source_sel == 14)) begin
        _tmp_464 <= read_rtl_bank_463;
      end 
      if(_stream_matmul_11_stream_oready && _stream_matmul_11_source_9_source_ram_renable && (_stream_matmul_11_source_9_source_sel == 2)) begin
        _tmp_1374 <= read_rtl_bank_1373;
      end 
    end
  end

  localparam _stream_conv2d_4_source_31_source_pat_fsm_13_1 = 1;
  localparam _stream_conv2d_4_source_31_source_pat_fsm_13_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_31_source_pat_fsm_13 <= _stream_conv2d_4_source_31_source_pat_fsm_13_init;
    end else begin
      case(_stream_conv2d_4_source_31_source_pat_fsm_13)
        _stream_conv2d_4_source_31_source_pat_fsm_13_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_31_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_31_source_pat_fsm_13 <= _stream_conv2d_4_source_31_source_pat_fsm_13_1;
          end 
        end
        _stream_conv2d_4_source_31_source_pat_fsm_13_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_31_source_pat_fsm_13 <= _stream_conv2d_4_source_31_source_pat_fsm_13_init;
          end 
          if((_source_stream_conv2d_4_source_31_pat_count_0 == 0) && (_source_stream_conv2d_4_source_31_pat_count_1 == 0) && (_source_stream_conv2d_4_source_31_pat_count_2 == 0) && (_source_stream_conv2d_4_source_31_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_31_source_pat_fsm_13 <= _stream_conv2d_4_source_31_source_pat_fsm_13_2;
          end 
        end
        _stream_conv2d_4_source_31_source_pat_fsm_13_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_31_source_pat_fsm_13 <= _stream_conv2d_4_source_31_source_pat_fsm_13_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_473 <= 0;
    end else begin
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_32_source_ram_renable && (_stream_conv2d_4_source_32_source_sel == 15)) begin
        _tmp_473 <= read_rtl_bank_472;
      end 
    end
  end

  localparam _stream_conv2d_4_source_32_source_pat_fsm_14_1 = 1;
  localparam _stream_conv2d_4_source_32_source_pat_fsm_14_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_32_source_pat_fsm_14 <= _stream_conv2d_4_source_32_source_pat_fsm_14_init;
    end else begin
      case(_stream_conv2d_4_source_32_source_pat_fsm_14)
        _stream_conv2d_4_source_32_source_pat_fsm_14_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_32_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_32_source_pat_fsm_14 <= _stream_conv2d_4_source_32_source_pat_fsm_14_1;
          end 
        end
        _stream_conv2d_4_source_32_source_pat_fsm_14_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_32_source_pat_fsm_14 <= _stream_conv2d_4_source_32_source_pat_fsm_14_init;
          end 
          if((_source_stream_conv2d_4_source_32_pat_count_0 == 0) && (_source_stream_conv2d_4_source_32_pat_count_1 == 0) && (_source_stream_conv2d_4_source_32_pat_count_2 == 0) && (_source_stream_conv2d_4_source_32_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_32_source_pat_fsm_14 <= _stream_conv2d_4_source_32_source_pat_fsm_14_2;
          end 
        end
        _stream_conv2d_4_source_32_source_pat_fsm_14_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_32_source_pat_fsm_14 <= _stream_conv2d_4_source_32_source_pat_fsm_14_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_482 <= 0;
    end else begin
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_33_source_ram_renable && (_stream_conv2d_4_source_33_source_sel == 16)) begin
        _tmp_482 <= read_rtl_bank_481;
      end 
    end
  end

  localparam _stream_conv2d_4_source_33_source_pat_fsm_15_1 = 1;
  localparam _stream_conv2d_4_source_33_source_pat_fsm_15_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_33_source_pat_fsm_15 <= _stream_conv2d_4_source_33_source_pat_fsm_15_init;
    end else begin
      case(_stream_conv2d_4_source_33_source_pat_fsm_15)
        _stream_conv2d_4_source_33_source_pat_fsm_15_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_33_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_33_source_pat_fsm_15 <= _stream_conv2d_4_source_33_source_pat_fsm_15_1;
          end 
        end
        _stream_conv2d_4_source_33_source_pat_fsm_15_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_33_source_pat_fsm_15 <= _stream_conv2d_4_source_33_source_pat_fsm_15_init;
          end 
          if((_source_stream_conv2d_4_source_33_pat_count_0 == 0) && (_source_stream_conv2d_4_source_33_pat_count_1 == 0) && (_source_stream_conv2d_4_source_33_pat_count_2 == 0) && (_source_stream_conv2d_4_source_33_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_33_source_pat_fsm_15 <= _stream_conv2d_4_source_33_source_pat_fsm_15_2;
          end 
        end
        _stream_conv2d_4_source_33_source_pat_fsm_15_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_33_source_pat_fsm_15 <= _stream_conv2d_4_source_33_source_pat_fsm_15_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_491 <= 0;
    end else begin
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_34_source_ram_renable && (_stream_conv2d_4_source_34_source_sel == 17)) begin
        _tmp_491 <= read_rtl_bank_490;
      end 
    end
  end

  localparam _stream_conv2d_4_source_34_source_pat_fsm_16_1 = 1;
  localparam _stream_conv2d_4_source_34_source_pat_fsm_16_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_34_source_pat_fsm_16 <= _stream_conv2d_4_source_34_source_pat_fsm_16_init;
    end else begin
      case(_stream_conv2d_4_source_34_source_pat_fsm_16)
        _stream_conv2d_4_source_34_source_pat_fsm_16_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_34_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_34_source_pat_fsm_16 <= _stream_conv2d_4_source_34_source_pat_fsm_16_1;
          end 
        end
        _stream_conv2d_4_source_34_source_pat_fsm_16_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_34_source_pat_fsm_16 <= _stream_conv2d_4_source_34_source_pat_fsm_16_init;
          end 
          if((_source_stream_conv2d_4_source_34_pat_count_0 == 0) && (_source_stream_conv2d_4_source_34_pat_count_1 == 0) && (_source_stream_conv2d_4_source_34_pat_count_2 == 0) && (_source_stream_conv2d_4_source_34_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_34_source_pat_fsm_16 <= _stream_conv2d_4_source_34_source_pat_fsm_16_2;
          end 
        end
        _stream_conv2d_4_source_34_source_pat_fsm_16_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_34_source_pat_fsm_16 <= _stream_conv2d_4_source_34_source_pat_fsm_16_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_500 <= 0;
    end else begin
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_35_source_ram_renable && (_stream_conv2d_4_source_35_source_sel == 18)) begin
        _tmp_500 <= read_rtl_bank_499;
      end 
    end
  end

  localparam _stream_conv2d_4_source_35_source_pat_fsm_17_1 = 1;
  localparam _stream_conv2d_4_source_35_source_pat_fsm_17_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_35_source_pat_fsm_17 <= _stream_conv2d_4_source_35_source_pat_fsm_17_init;
    end else begin
      case(_stream_conv2d_4_source_35_source_pat_fsm_17)
        _stream_conv2d_4_source_35_source_pat_fsm_17_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_35_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_35_source_pat_fsm_17 <= _stream_conv2d_4_source_35_source_pat_fsm_17_1;
          end 
        end
        _stream_conv2d_4_source_35_source_pat_fsm_17_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_35_source_pat_fsm_17 <= _stream_conv2d_4_source_35_source_pat_fsm_17_init;
          end 
          if((_source_stream_conv2d_4_source_35_pat_count_0 == 0) && (_source_stream_conv2d_4_source_35_pat_count_1 == 0) && (_source_stream_conv2d_4_source_35_pat_count_2 == 0) && (_source_stream_conv2d_4_source_35_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_35_source_pat_fsm_17 <= _stream_conv2d_4_source_35_source_pat_fsm_17_2;
          end 
        end
        _stream_conv2d_4_source_35_source_pat_fsm_17_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_35_source_pat_fsm_17 <= _stream_conv2d_4_source_35_source_pat_fsm_17_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_509 <= 0;
    end else begin
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_36_source_ram_renable && (_stream_conv2d_4_source_36_source_sel == 19)) begin
        _tmp_509 <= read_rtl_bank_508;
      end 
    end
  end

  localparam _stream_conv2d_4_source_36_source_pat_fsm_18_1 = 1;
  localparam _stream_conv2d_4_source_36_source_pat_fsm_18_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_36_source_pat_fsm_18 <= _stream_conv2d_4_source_36_source_pat_fsm_18_init;
    end else begin
      case(_stream_conv2d_4_source_36_source_pat_fsm_18)
        _stream_conv2d_4_source_36_source_pat_fsm_18_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_36_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_36_source_pat_fsm_18 <= _stream_conv2d_4_source_36_source_pat_fsm_18_1;
          end 
        end
        _stream_conv2d_4_source_36_source_pat_fsm_18_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_36_source_pat_fsm_18 <= _stream_conv2d_4_source_36_source_pat_fsm_18_init;
          end 
          if((_source_stream_conv2d_4_source_36_pat_count_0 == 0) && (_source_stream_conv2d_4_source_36_pat_count_1 == 0) && (_source_stream_conv2d_4_source_36_pat_count_2 == 0) && (_source_stream_conv2d_4_source_36_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_36_source_pat_fsm_18 <= _stream_conv2d_4_source_36_source_pat_fsm_18_2;
          end 
        end
        _stream_conv2d_4_source_36_source_pat_fsm_18_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_36_source_pat_fsm_18 <= _stream_conv2d_4_source_36_source_pat_fsm_18_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_518 <= 0;
    end else begin
      if(_stream_conv2d_4_stream_oready && _stream_conv2d_4_source_37_source_ram_renable && (_stream_conv2d_4_source_37_source_sel == 20)) begin
        _tmp_518 <= read_rtl_bank_517;
      end 
    end
  end

  localparam _stream_conv2d_4_source_37_source_pat_fsm_19_1 = 1;
  localparam _stream_conv2d_4_source_37_source_pat_fsm_19_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_source_37_source_pat_fsm_19 <= _stream_conv2d_4_source_37_source_pat_fsm_19_init;
    end else begin
      case(_stream_conv2d_4_source_37_source_pat_fsm_19)
        _stream_conv2d_4_source_37_source_pat_fsm_19_init: begin
          if(_stream_conv2d_4_source_start && _stream_conv2d_4_source_37_source_mode & 5'b10 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_37_source_pat_fsm_19 <= _stream_conv2d_4_source_37_source_pat_fsm_19_1;
          end 
        end
        _stream_conv2d_4_source_37_source_pat_fsm_19_1: begin
          if(_stream_conv2d_4_source_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_37_source_pat_fsm_19 <= _stream_conv2d_4_source_37_source_pat_fsm_19_init;
          end 
          if((_source_stream_conv2d_4_source_37_pat_count_0 == 0) && (_source_stream_conv2d_4_source_37_pat_count_1 == 0) && (_source_stream_conv2d_4_source_37_pat_count_2 == 0) && (_source_stream_conv2d_4_source_37_pat_count_3 == 0) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_37_source_pat_fsm_19 <= _stream_conv2d_4_source_37_source_pat_fsm_19_2;
          end 
        end
        _stream_conv2d_4_source_37_source_pat_fsm_19_2: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_source_37_source_pat_fsm_19 <= _stream_conv2d_4_source_37_source_pat_fsm_19_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_conv2d_4_sink_50_sink_fsm_20_1 = 1;
  localparam _stream_conv2d_4_sink_50_sink_fsm_20_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_conv2d_4_sink_50_sink_fsm_20 <= _stream_conv2d_4_sink_50_sink_fsm_20_init;
    end else begin
      case(_stream_conv2d_4_sink_50_sink_fsm_20)
        _stream_conv2d_4_sink_50_sink_fsm_20_init: begin
          if(_stream_conv2d_4_sink_start && _stream_conv2d_4_sink_50_sink_mode & 5'b1 && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_sink_50_sink_fsm_20 <= _stream_conv2d_4_sink_50_sink_fsm_20_1;
          end 
        end
        _stream_conv2d_4_sink_50_sink_fsm_20_1: begin
          if(_stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_sink_50_sink_fsm_20 <= _stream_conv2d_4_sink_50_sink_fsm_20_2;
          end 
        end
        _stream_conv2d_4_sink_50_sink_fsm_20_2: begin
          if(stream_conv2d_4_sink_51_data && (_stream_conv2d_4_sink_50_sink_count == 1) && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_sink_50_sink_fsm_20 <= _stream_conv2d_4_sink_50_sink_fsm_20_init;
          end 
          if(_stream_conv2d_4_sink_stop && _stream_conv2d_4_stream_oready) begin
            _stream_conv2d_4_sink_50_sink_fsm_20 <= _stream_conv2d_4_sink_50_sink_fsm_20_init;
          end 
        end
      endcase
    end
  end

  localparam _maxi_write_req_fsm_1 = 1;

  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _maxi_write_req_fsm <= _maxi_write_req_fsm_init;
      _maxi_write_cont <= 0;
    end else begin
      case(_maxi_write_req_fsm)
        _maxi_write_req_fsm_init: begin
          if((_maxi_write_req_fsm == 0) && (_maxi_write_start || _maxi_write_cont) && !_maxi_write_req_fifo_almost_full) begin
            _maxi_write_req_fsm <= _maxi_write_req_fsm_1;
          end 
        end
        _maxi_write_req_fsm_1: begin
          if((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (maxi_awready || !maxi_awvalid) && (_maxi_outstanding_wcount < 6)) begin
            _maxi_write_cont <= 1;
          end 
          if((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (maxi_awready || !maxi_awvalid) && (_maxi_outstanding_wcount < 6) && (_maxi_write_global_size == 0)) begin
            _maxi_write_cont <= 0;
          end 
          if((_maxi_write_req_fsm == 1) && !_maxi_write_req_fifo_almost_full && (maxi_awready || !maxi_awvalid) && (_maxi_outstanding_wcount < 6)) begin
            _maxi_write_req_fsm <= _maxi_write_req_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam _maxi_write_data_fsm_1 = 1;
  localparam _maxi_write_data_fsm_2 = 2;

  always @(posedge CLK) begin
    if(RESETN_inv_buf) begin
      _maxi_write_data_fsm <= _maxi_write_data_fsm_init;
    end else begin
      case(_maxi_write_data_fsm)
        _maxi_write_data_fsm_init: begin
          if(!_maxi_write_data_busy && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 1)) begin
            _maxi_write_data_fsm <= _maxi_write_data_fsm_1;
          end 
          if(!_maxi_write_data_busy && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 2)) begin
            _maxi_write_data_fsm <= _maxi_write_data_fsm_1;
          end 
          if(!_maxi_write_data_busy && !_maxi_write_req_fifo_empty && (_maxi_write_op_sel_fifo == 3)) begin
            _maxi_write_data_fsm <= _maxi_write_data_fsm_1;
          end 
        end
        _maxi_write_data_fsm_1: begin
          _maxi_write_data_fsm <= _maxi_write_data_fsm_2;
          _maxi_write_data_fsm <= _maxi_write_data_fsm_2;
          _maxi_write_data_fsm <= _maxi_write_data_fsm_2;
        end
        _maxi_write_data_fsm_2: begin
          if((_maxi_write_op_sel_buf == 1) && read_burst_packed_rvalid_1169 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)) && read_burst_packed_rlast_1170) begin
            _maxi_write_data_fsm <= _maxi_write_data_fsm_init;
          end 
          if((_maxi_write_op_sel_buf == 2) && read_burst_packed_rvalid_1301 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)) && read_burst_packed_rlast_1302) begin
            _maxi_write_data_fsm <= _maxi_write_data_fsm_init;
          end 
          if((_maxi_write_op_sel_buf == 3) && read_burst_packed_rvalid_1635 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0)) && read_burst_packed_rlast_1636) begin
            _maxi_write_data_fsm <= _maxi_write_data_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam read_burst_packed_fsm_55_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      read_burst_packed_fsm_55 <= read_burst_packed_fsm_55_init;
      read_burst_packed_addr_1166 <= 0;
      read_burst_packed_stride_1167 <= 0;
      read_burst_packed_length_1168 <= 0;
      read_burst_packed_rvalid_1169 <= 0;
      read_burst_packed_rlast_1170 <= 0;
    end else begin
      case(read_burst_packed_fsm_55)
        read_burst_packed_fsm_55_init: begin
          read_burst_packed_addr_1166 <= _maxi_write_local_addr_buf;
          read_burst_packed_stride_1167 <= _maxi_write_local_stride_buf;
          read_burst_packed_length_1168 <= _maxi_write_size_buf;
          read_burst_packed_rvalid_1169 <= 0;
          read_burst_packed_rlast_1170 <= 0;
          if((_maxi_write_data_fsm == 1) && (_maxi_write_op_sel_buf == 1) && (_maxi_write_size_buf > 0)) begin
            read_burst_packed_fsm_55 <= read_burst_packed_fsm_55_1;
          end 
        end
        read_burst_packed_fsm_55_1: begin
          if((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0) && (read_burst_packed_length_1168 > 0)) begin
            read_burst_packed_addr_1166 <= read_burst_packed_addr_1166 + read_burst_packed_stride_1167;
            read_burst_packed_length_1168 <= read_burst_packed_length_1168 - 1;
            read_burst_packed_rvalid_1169 <= 1;
          end 
          if((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0) && (read_burst_packed_length_1168 <= 1)) begin
            read_burst_packed_rlast_1170 <= 1;
          end 
          if(read_burst_packed_rlast_1170 && read_burst_packed_rvalid_1169 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) begin
            read_burst_packed_rvalid_1169 <= 0;
            read_burst_packed_rlast_1170 <= 0;
          end 
          if(0) begin
            read_burst_packed_rvalid_1169 <= 0;
            read_burst_packed_rlast_1170 <= 0;
          end 
          if(read_burst_packed_rlast_1170 && read_burst_packed_rvalid_1169 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) begin
            read_burst_packed_fsm_55 <= read_burst_packed_fsm_55_init;
          end 
          if(0) begin
            read_burst_packed_fsm_55 <= read_burst_packed_fsm_55_init;
          end 
        end
      endcase
    end
  end

  localparam control_max_pool_serial_6_1 = 1;
  localparam control_max_pool_serial_6_2 = 2;
  localparam control_max_pool_serial_6_3 = 3;
  localparam control_max_pool_serial_6_4 = 4;
  localparam control_max_pool_serial_6_5 = 5;
  localparam control_max_pool_serial_6_6 = 6;
  localparam control_max_pool_serial_6_7 = 7;
  localparam control_max_pool_serial_6_8 = 8;
  localparam control_max_pool_serial_6_9 = 9;
  localparam control_max_pool_serial_6_10 = 10;
  localparam control_max_pool_serial_6_11 = 11;
  localparam control_max_pool_serial_6_12 = 12;
  localparam control_max_pool_serial_6_13 = 13;
  localparam control_max_pool_serial_6_14 = 14;
  localparam control_max_pool_serial_6_15 = 15;
  localparam control_max_pool_serial_6_16 = 16;
  localparam control_max_pool_serial_6_17 = 17;
  localparam control_max_pool_serial_6_18 = 18;
  localparam control_max_pool_serial_6_19 = 19;

  always @(posedge CLK) begin
    if(RST) begin
      control_max_pool_serial_6 <= control_max_pool_serial_6_init;
      _control_max_pool_serial_6_called <= 0;
      max_pool_serial_6_act_base_offset_row <= 0;
      max_pool_serial_6_act_base_offset_bat <= 0;
      max_pool_serial_6_act_page <= 0;
      max_pool_serial_6_act_page_comp_offset <= 0;
      max_pool_serial_6_act_page_dma_offset <= 0;
      max_pool_serial_6_out_base_offset_row <= 0;
      max_pool_serial_6_out_base_offset_bat <= 0;
      max_pool_serial_6_out_page <= 0;
      max_pool_serial_6_out_page_comp_offset <= 0;
      max_pool_serial_6_out_page_dma_offset <= 0;
      max_pool_serial_6_row_count <= 0;
      max_pool_serial_6_bat_count <= 0;
      max_pool_serial_6_prev_row_count <= 0;
      max_pool_serial_6_prev_bat_count <= 0;
      max_pool_serial_6_skip_read_act <= 0;
      max_pool_serial_6_skip_comp <= 0;
      max_pool_serial_6_skip_write_out <= 0;
      max_pool_serial_6_out_count <= 0;
    end else begin
      case(control_max_pool_serial_6)
        control_max_pool_serial_6_init: begin
          if(main_fsm == 16) begin
            _control_max_pool_serial_6_called <= 1;
          end 
          if(main_fsm == 16) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_1;
          end 
        end
        control_max_pool_serial_6_1: begin
          control_max_pool_serial_6 <= control_max_pool_serial_6_2;
        end
        control_max_pool_serial_6_2: begin
          max_pool_serial_6_act_base_offset_row <= 0;
          max_pool_serial_6_act_base_offset_bat <= 0;
          max_pool_serial_6_act_page <= 0;
          max_pool_serial_6_act_page_comp_offset <= 0;
          max_pool_serial_6_act_page_dma_offset <= 0;
          max_pool_serial_6_out_base_offset_row <= 0;
          max_pool_serial_6_out_base_offset_bat <= 0;
          max_pool_serial_6_out_page <= 0;
          max_pool_serial_6_out_page_comp_offset <= 0;
          max_pool_serial_6_out_page_dma_offset <= 0;
          max_pool_serial_6_row_count <= 0;
          max_pool_serial_6_bat_count <= 0;
          max_pool_serial_6_prev_row_count <= 0;
          max_pool_serial_6_prev_bat_count <= 0;
          max_pool_serial_6_skip_read_act <= 0;
          max_pool_serial_6_skip_comp <= 0;
          max_pool_serial_6_skip_write_out <= 1;
          max_pool_serial_6_out_count <= 0;
          control_max_pool_serial_6 <= control_max_pool_serial_6_3;
        end
        control_max_pool_serial_6_3: begin
          control_max_pool_serial_6 <= control_max_pool_serial_6_4;
          if(max_pool_serial_6_skip_read_act) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_11;
          end 
        end
        control_max_pool_serial_6_4: begin
          control_max_pool_serial_6 <= control_max_pool_serial_6_5;
          if(max_pool_serial_6_dma_pad_mask_0) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_7;
          end 
        end
        control_max_pool_serial_6_5: begin
          if(_maxi_read_req_idle) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_6;
          end 
        end
        control_max_pool_serial_6_6: begin
          if(_maxi_read_idle) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_7;
          end 
        end
        control_max_pool_serial_6_7: begin
          control_max_pool_serial_6 <= control_max_pool_serial_6_8;
          if(max_pool_serial_6_dma_pad_mask_1) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_10;
          end 
        end
        control_max_pool_serial_6_8: begin
          if(_maxi_read_req_idle) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_9;
          end 
        end
        control_max_pool_serial_6_9: begin
          if(_maxi_read_idle) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_10;
          end 
        end
        control_max_pool_serial_6_10: begin
          control_max_pool_serial_6 <= control_max_pool_serial_6_11;
        end
        control_max_pool_serial_6_11: begin
          if(_maxi_write_idle) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_12;
          end 
        end
        control_max_pool_serial_6_12: begin
          if(max_pool_serial_6_comp_fsm == 0) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_13;
          end 
        end
        control_max_pool_serial_6_13: begin
          control_max_pool_serial_6 <= control_max_pool_serial_6_14;
          if(max_pool_serial_6_skip_write_out) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_17;
          end 
        end
        control_max_pool_serial_6_14: begin
          if(max_pool_serial_6_comp_count >= max_pool_serial_6_out_count + cparam_max_pool_serial_6_out_write_size) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_15;
          end 
        end
        control_max_pool_serial_6_15: begin
          if(_maxi_write_req_idle) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_16;
          end 
        end
        control_max_pool_serial_6_16: begin
          max_pool_serial_6_out_count <= max_pool_serial_6_out_count + cparam_max_pool_serial_6_out_write_size;
          control_max_pool_serial_6 <= control_max_pool_serial_6_17;
        end
        control_max_pool_serial_6_17: begin
          max_pool_serial_6_act_base_offset_row <= max_pool_serial_6_act_base_offset_row + cparam_max_pool_serial_6_act_row_step;
          if(max_pool_serial_6_row_count >= cparam_max_pool_serial_6_max_row_count) begin
            max_pool_serial_6_act_base_offset_row <= 0;
            max_pool_serial_6_act_base_offset_bat <= max_pool_serial_6_act_base_offset_bat + cparam_max_pool_serial_6_act_bat_step;
          end 
          if((max_pool_serial_6_row_count >= cparam_max_pool_serial_6_max_row_count) && (max_pool_serial_6_bat_count >= cparam_max_pool_serial_6_max_bat_count)) begin
            max_pool_serial_6_act_base_offset_bat <= 0;
          end 
          max_pool_serial_6_row_count <= max_pool_serial_6_row_count + cparam_max_pool_serial_6_stride_row;
          if(max_pool_serial_6_row_count >= cparam_max_pool_serial_6_max_row_count) begin
            max_pool_serial_6_row_count <= 0;
            max_pool_serial_6_bat_count <= max_pool_serial_6_bat_count + 1;
          end 
          if((max_pool_serial_6_row_count >= cparam_max_pool_serial_6_max_row_count) && (max_pool_serial_6_bat_count >= cparam_max_pool_serial_6_max_bat_count)) begin
            max_pool_serial_6_bat_count <= 0;
          end 
          if(!max_pool_serial_6_act_page) begin
            max_pool_serial_6_act_page_comp_offset <= 16384;
            max_pool_serial_6_act_page_dma_offset <= 16384;
            max_pool_serial_6_act_page <= 1;
          end 
          if(max_pool_serial_6_act_page) begin
            max_pool_serial_6_act_page_comp_offset <= 0;
            max_pool_serial_6_act_page_dma_offset <= 0;
            max_pool_serial_6_act_page <= 0;
          end 
          if(!max_pool_serial_6_skip_write_out) begin
            max_pool_serial_6_out_base_offset_row <= max_pool_serial_6_out_base_offset_row + cparam_max_pool_serial_6_out_row_step;
          end 
          if(!max_pool_serial_6_skip_write_out && (max_pool_serial_6_prev_row_count >= cparam_max_pool_serial_6_max_row_count)) begin
            max_pool_serial_6_out_base_offset_row <= 0;
            max_pool_serial_6_out_base_offset_bat <= max_pool_serial_6_out_base_offset_bat + cparam_max_pool_serial_6_out_bat_step;
          end 
          if(!max_pool_serial_6_skip_write_out && (max_pool_serial_6_prev_row_count >= cparam_max_pool_serial_6_max_row_count) && (max_pool_serial_6_prev_bat_count >= cparam_max_pool_serial_6_max_bat_count)) begin
            max_pool_serial_6_out_base_offset_bat <= 0;
          end 
          if(!max_pool_serial_6_out_page) begin
            max_pool_serial_6_out_page_comp_offset <= 4096;
            max_pool_serial_6_out_page_dma_offset <= 0;
            max_pool_serial_6_out_page <= 1;
          end 
          if(max_pool_serial_6_out_page) begin
            max_pool_serial_6_out_page_comp_offset <= 0;
            max_pool_serial_6_out_page_dma_offset <= 4096;
            max_pool_serial_6_out_page <= 0;
          end 
          max_pool_serial_6_prev_row_count <= max_pool_serial_6_row_count;
          max_pool_serial_6_prev_bat_count <= max_pool_serial_6_bat_count;
          if((max_pool_serial_6_row_count >= cparam_max_pool_serial_6_max_row_count) && (max_pool_serial_6_bat_count >= cparam_max_pool_serial_6_max_bat_count)) begin
            max_pool_serial_6_skip_read_act <= 1;
          end 
          if((max_pool_serial_6_row_count >= cparam_max_pool_serial_6_max_row_count) && (max_pool_serial_6_bat_count >= cparam_max_pool_serial_6_max_bat_count)) begin
            max_pool_serial_6_skip_comp <= 1;
          end 
          if(max_pool_serial_6_skip_write_out && (max_pool_serial_6_prev_row_count == 0) && (max_pool_serial_6_prev_bat_count == 0)) begin
            max_pool_serial_6_skip_write_out <= 0;
          end 
          control_max_pool_serial_6 <= control_max_pool_serial_6_3;
          if(!max_pool_serial_6_skip_write_out && (max_pool_serial_6_prev_row_count >= cparam_max_pool_serial_6_max_row_count) && (max_pool_serial_6_prev_bat_count >= cparam_max_pool_serial_6_max_bat_count)) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_18;
          end 
        end
        control_max_pool_serial_6_18: begin
          if(_maxi_write_idle && !_maxi_has_outstanding_write) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_19;
          end 
        end
        control_max_pool_serial_6_19: begin
          if(main_fsm == 19) begin
            _control_max_pool_serial_6_called <= 0;
          end 
          if(main_fsm == 19) begin
            control_max_pool_serial_6 <= control_max_pool_serial_6_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_56_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_56 <= write_burst_packed_fsm_56_init;
      write_burst_packed_addr_1185 <= 0;
      write_burst_packed_stride_1186 <= 0;
      write_burst_packed_length_1187 <= 0;
      write_burst_packed_done_1188 <= 0;
    end else begin
      case(write_burst_packed_fsm_56)
        write_burst_packed_fsm_56_init: begin
          write_burst_packed_addr_1185 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_1186 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_1187 <= _maxi_read_local_size_buf;
          write_burst_packed_done_1188 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 7) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_56 <= write_burst_packed_fsm_56_1;
          end 
        end
        write_burst_packed_fsm_56_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_packed_addr_1185 <= write_burst_packed_addr_1185 + write_burst_packed_stride_1186;
            write_burst_packed_length_1187 <= write_burst_packed_length_1187 - 1;
            write_burst_packed_done_1188 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_packed_length_1187 <= 1)) begin
            write_burst_packed_done_1188 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_packed_done_1188 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_packed_length_1187 <= 1)) begin
            write_burst_packed_fsm_56 <= write_burst_packed_fsm_56_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_packed_fsm_56 <= write_burst_packed_fsm_56_init;
          end 
          if(0) begin
            write_burst_packed_fsm_56 <= write_burst_packed_fsm_56_init;
          end 
        end
      endcase
    end
  end

  localparam max_pool_serial_6_comp_fsm_1 = 1;
  localparam max_pool_serial_6_comp_fsm_2 = 2;
  localparam max_pool_serial_6_comp_fsm_3 = 3;
  localparam max_pool_serial_6_comp_fsm_4 = 4;
  localparam max_pool_serial_6_comp_fsm_5 = 5;
  localparam max_pool_serial_6_comp_fsm_6 = 6;
  localparam max_pool_serial_6_comp_fsm_7 = 7;

  always @(posedge CLK) begin
    if(RST) begin
      max_pool_serial_6_comp_fsm <= max_pool_serial_6_comp_fsm_init;
      max_pool_serial_6_stream_act_local <= 0;
      max_pool_serial_6_stream_out_local <= 0;
      max_pool_serial_6_col_count <= 0;
      max_pool_serial_6_act_page_comp_offset_buf <= 0;
      max_pool_serial_6_out_page_comp_offset_buf <= 0;
      max_pool_serial_6_row_count_buf <= 0;
      max_pool_serial_6_stream_pad_masks <= 0;
      max_pool_serial_6_comp_count <= 0;
    end else begin
      if(control_max_pool_serial_6 == 2) begin
        max_pool_serial_6_comp_count <= 0;
      end 
      if(_stream_max_pool_serial_6_sink_stop) begin
        max_pool_serial_6_comp_count <= max_pool_serial_6_comp_count + cparam_max_pool_serial_6_inc_out_laddr;
      end 
      case(max_pool_serial_6_comp_fsm)
        max_pool_serial_6_comp_fsm_init: begin
          if((control_max_pool_serial_6 == 12) && !max_pool_serial_6_skip_comp) begin
            max_pool_serial_6_comp_fsm <= max_pool_serial_6_comp_fsm_1;
          end 
        end
        max_pool_serial_6_comp_fsm_1: begin
          max_pool_serial_6_stream_act_local <= cparam_max_pool_serial_6_local_pad_offset;
          max_pool_serial_6_stream_out_local <= 0;
          max_pool_serial_6_col_count <= 0;
          max_pool_serial_6_act_page_comp_offset_buf <= max_pool_serial_6_act_page_comp_offset;
          max_pool_serial_6_out_page_comp_offset_buf <= max_pool_serial_6_out_page_comp_offset;
          max_pool_serial_6_row_count_buf <= max_pool_serial_6_row_count;
          max_pool_serial_6_comp_fsm <= max_pool_serial_6_comp_fsm_2;
        end
        max_pool_serial_6_comp_fsm_2: begin
          max_pool_serial_6_stream_pad_masks <= { max_pool_serial_6_stream_pad_mask_1_1, max_pool_serial_6_stream_pad_mask_1_0, max_pool_serial_6_stream_pad_mask_0_1, max_pool_serial_6_stream_pad_mask_0_0 };
          max_pool_serial_6_comp_fsm <= max_pool_serial_6_comp_fsm_3;
        end
        max_pool_serial_6_comp_fsm_3: begin
          if(!_stream_max_pool_serial_6_source_busy) begin
            max_pool_serial_6_comp_fsm <= max_pool_serial_6_comp_fsm_4;
          end 
        end
        max_pool_serial_6_comp_fsm_4: begin
          max_pool_serial_6_comp_fsm <= max_pool_serial_6_comp_fsm_5;
          max_pool_serial_6_comp_fsm <= max_pool_serial_6_comp_fsm_5;
          max_pool_serial_6_comp_fsm <= max_pool_serial_6_comp_fsm_5;
          if(_stream_max_pool_serial_6_stream_oready) begin
            max_pool_serial_6_comp_fsm <= max_pool_serial_6_comp_fsm_5;
          end 
        end
        max_pool_serial_6_comp_fsm_5: begin
          max_pool_serial_6_comp_fsm <= max_pool_serial_6_comp_fsm_6;
        end
        max_pool_serial_6_comp_fsm_6: begin
          if(_stream_max_pool_serial_6_busy) begin
            max_pool_serial_6_comp_fsm <= max_pool_serial_6_comp_fsm_7;
          end 
        end
        max_pool_serial_6_comp_fsm_7: begin
          max_pool_serial_6_stream_act_local <= max_pool_serial_6_stream_act_local + cparam_max_pool_serial_6_inc_act_laddr;
          if(max_pool_serial_6_col_count >= cparam_max_pool_serial_6_max_col_count) begin
            max_pool_serial_6_stream_act_local <= cparam_max_pool_serial_6_local_pad_offset;
          end 
          max_pool_serial_6_stream_out_local <= max_pool_serial_6_stream_out_local + cparam_max_pool_serial_6_inc_out_laddr;
          if(max_pool_serial_6_col_count >= cparam_max_pool_serial_6_max_col_count) begin
            max_pool_serial_6_stream_out_local <= 0;
          end 
          max_pool_serial_6_col_count <= max_pool_serial_6_col_count + cparam_max_pool_serial_6_stride_col;
          if(max_pool_serial_6_col_count >= cparam_max_pool_serial_6_max_col_count) begin
            max_pool_serial_6_col_count <= 0;
          end 
          max_pool_serial_6_comp_fsm <= max_pool_serial_6_comp_fsm_2;
          if(max_pool_serial_6_col_count >= cparam_max_pool_serial_6_max_col_count) begin
            max_pool_serial_6_comp_fsm <= max_pool_serial_6_comp_fsm_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_1202 <= 0;
      _tmp_1402 <= 0;
    end else begin
      if(_stream_max_pool_serial_6_stream_oready && _stream_max_pool_serial_6_source_1_source_ram_renable && (_stream_max_pool_serial_6_source_1_source_sel == 1)) begin
        _tmp_1202 <= read_rtl_bank_1201;
      end 
      if(_stream_matmul_11_stream_oready && _stream_matmul_11_source_21_source_ram_renable && (_stream_matmul_11_source_21_source_sel == 4)) begin
        _tmp_1402 <= read_rtl_bank_1401;
      end 
    end
  end

  localparam _stream_max_pool_serial_6_source_1_source_pat_fsm_0_1 = 1;
  localparam _stream_max_pool_serial_6_source_1_source_pat_fsm_0_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_max_pool_serial_6_source_1_source_pat_fsm_0 <= _stream_max_pool_serial_6_source_1_source_pat_fsm_0_init;
    end else begin
      case(_stream_max_pool_serial_6_source_1_source_pat_fsm_0)
        _stream_max_pool_serial_6_source_1_source_pat_fsm_0_init: begin
          if(_stream_max_pool_serial_6_source_start && _stream_max_pool_serial_6_source_1_source_mode & 5'b10 && _stream_max_pool_serial_6_stream_oready) begin
            _stream_max_pool_serial_6_source_1_source_pat_fsm_0 <= _stream_max_pool_serial_6_source_1_source_pat_fsm_0_1;
          end 
        end
        _stream_max_pool_serial_6_source_1_source_pat_fsm_0_1: begin
          if(_stream_max_pool_serial_6_source_stop && _stream_max_pool_serial_6_stream_oready) begin
            _stream_max_pool_serial_6_source_1_source_pat_fsm_0 <= _stream_max_pool_serial_6_source_1_source_pat_fsm_0_init;
          end 
          if((_source_stream_max_pool_serial_6_source_1_pat_count_0 == 0) && (_source_stream_max_pool_serial_6_source_1_pat_count_1 == 0) && (_source_stream_max_pool_serial_6_source_1_pat_count_2 == 0) && (_source_stream_max_pool_serial_6_source_1_pat_count_3 == 0) && _stream_max_pool_serial_6_stream_oready) begin
            _stream_max_pool_serial_6_source_1_source_pat_fsm_0 <= _stream_max_pool_serial_6_source_1_source_pat_fsm_0_2;
          end 
        end
        _stream_max_pool_serial_6_source_1_source_pat_fsm_0_2: begin
          if(_stream_max_pool_serial_6_stream_oready) begin
            _stream_max_pool_serial_6_source_1_source_pat_fsm_0 <= _stream_max_pool_serial_6_source_1_source_pat_fsm_0_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_max_pool_serial_6_sink_5_sink_fsm_1_1 = 1;
  localparam _stream_max_pool_serial_6_sink_5_sink_fsm_1_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_max_pool_serial_6_sink_5_sink_fsm_1 <= _stream_max_pool_serial_6_sink_5_sink_fsm_1_init;
    end else begin
      case(_stream_max_pool_serial_6_sink_5_sink_fsm_1)
        _stream_max_pool_serial_6_sink_5_sink_fsm_1_init: begin
          if(_stream_max_pool_serial_6_sink_start && _stream_max_pool_serial_6_sink_5_sink_mode & 5'b1 && _stream_max_pool_serial_6_stream_oready) begin
            _stream_max_pool_serial_6_sink_5_sink_fsm_1 <= _stream_max_pool_serial_6_sink_5_sink_fsm_1_1;
          end 
        end
        _stream_max_pool_serial_6_sink_5_sink_fsm_1_1: begin
          if(_stream_max_pool_serial_6_stream_oready) begin
            _stream_max_pool_serial_6_sink_5_sink_fsm_1 <= _stream_max_pool_serial_6_sink_5_sink_fsm_1_2;
          end 
        end
        _stream_max_pool_serial_6_sink_5_sink_fsm_1_2: begin
          if(stream_max_pool_serial_6_sink_6_data && (_stream_max_pool_serial_6_sink_5_sink_count == 1) && _stream_max_pool_serial_6_stream_oready) begin
            _stream_max_pool_serial_6_sink_5_sink_fsm_1 <= _stream_max_pool_serial_6_sink_5_sink_fsm_1_init;
          end 
          if(_stream_max_pool_serial_6_sink_stop && _stream_max_pool_serial_6_stream_oready) begin
            _stream_max_pool_serial_6_sink_5_sink_fsm_1 <= _stream_max_pool_serial_6_sink_5_sink_fsm_1_init;
          end 
        end
      endcase
    end
  end

  localparam read_burst_packed_fsm_57_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      read_burst_packed_fsm_57 <= read_burst_packed_fsm_57_init;
      read_burst_packed_addr_1298 <= 0;
      read_burst_packed_stride_1299 <= 0;
      read_burst_packed_length_1300 <= 0;
      read_burst_packed_rvalid_1301 <= 0;
      read_burst_packed_rlast_1302 <= 0;
    end else begin
      case(read_burst_packed_fsm_57)
        read_burst_packed_fsm_57_init: begin
          read_burst_packed_addr_1298 <= _maxi_write_local_addr_buf;
          read_burst_packed_stride_1299 <= _maxi_write_local_stride_buf;
          read_burst_packed_length_1300 <= _maxi_write_size_buf;
          read_burst_packed_rvalid_1301 <= 0;
          read_burst_packed_rlast_1302 <= 0;
          if((_maxi_write_data_fsm == 1) && (_maxi_write_op_sel_buf == 2) && (_maxi_write_size_buf > 0)) begin
            read_burst_packed_fsm_57 <= read_burst_packed_fsm_57_1;
          end 
        end
        read_burst_packed_fsm_57_1: begin
          if((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0) && (read_burst_packed_length_1300 > 0)) begin
            read_burst_packed_addr_1298 <= read_burst_packed_addr_1298 + read_burst_packed_stride_1299;
            read_burst_packed_length_1300 <= read_burst_packed_length_1300 - 1;
            read_burst_packed_rvalid_1301 <= 1;
          end 
          if((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0) && (read_burst_packed_length_1300 <= 1)) begin
            read_burst_packed_rlast_1302 <= 1;
          end 
          if(read_burst_packed_rlast_1302 && read_burst_packed_rvalid_1301 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) begin
            read_burst_packed_rvalid_1301 <= 0;
            read_burst_packed_rlast_1302 <= 0;
          end 
          if(0) begin
            read_burst_packed_rvalid_1301 <= 0;
            read_burst_packed_rlast_1302 <= 0;
          end 
          if(read_burst_packed_rlast_1302 && read_burst_packed_rvalid_1301 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) begin
            read_burst_packed_fsm_57 <= read_burst_packed_fsm_57_init;
          end 
          if(0) begin
            read_burst_packed_fsm_57 <= read_burst_packed_fsm_57_init;
          end 
        end
      endcase
    end
  end

  localparam control_matmul_11_1 = 1;
  localparam control_matmul_11_2 = 2;
  localparam control_matmul_11_3 = 3;
  localparam control_matmul_11_4 = 4;
  localparam control_matmul_11_5 = 5;
  localparam control_matmul_11_6 = 6;
  localparam control_matmul_11_7 = 7;
  localparam control_matmul_11_8 = 8;
  localparam control_matmul_11_9 = 9;
  localparam control_matmul_11_10 = 10;
  localparam control_matmul_11_11 = 11;
  localparam control_matmul_11_12 = 12;
  localparam control_matmul_11_13 = 13;
  localparam control_matmul_11_14 = 14;
  localparam control_matmul_11_15 = 15;
  localparam control_matmul_11_16 = 16;
  localparam control_matmul_11_17 = 17;
  localparam control_matmul_11_18 = 18;
  localparam control_matmul_11_19 = 19;
  localparam control_matmul_11_20 = 20;
  localparam control_matmul_11_21 = 21;
  localparam control_matmul_11_22 = 22;
  localparam control_matmul_11_23 = 23;
  localparam control_matmul_11_24 = 24;
  localparam control_matmul_11_25 = 25;
  localparam control_matmul_11_26 = 26;
  localparam control_matmul_11_27 = 27;
  localparam control_matmul_11_28 = 28;

  always @(posedge CLK) begin
    if(RST) begin
      control_matmul_11 <= control_matmul_11_init;
      _control_matmul_11_called <= 0;
      matmul_11_filter_base_offset <= 0;
      matmul_11_filter_page_comp_offset <= 0;
      matmul_11_filter_page_dma_offset <= 0;
      matmul_11_act_base_offset_row <= 0;
      matmul_11_act_base_offset_bat <= 0;
      matmul_11_dma_flag_0 <= 0;
      matmul_11_act_page_comp_offset_0 <= 0;
      matmul_11_act_page_dma_offset_0 <= 0;
      matmul_11_out_base_offset_val <= 0;
      matmul_11_out_base_offset_col <= 0;
      matmul_11_out_base_offset_row <= 0;
      matmul_11_out_base_offset_bat <= 0;
      matmul_11_out_base_offset_och <= 0;
      matmul_11_out_page <= 0;
      matmul_11_out_page_comp_offset <= 0;
      matmul_11_out_page_dma_offset <= 0;
      matmul_11_out_laddr_offset <= 0;
      matmul_11_sync_out_count <= 0;
      matmul_11_write_count <= 0;
      matmul_11_next_out_write_size <= 0;
      matmul_11_row_count <= 0;
      matmul_11_bat_count <= 0;
      matmul_11_och_count <= 0;
      matmul_11_row_select <= 0;
      matmul_11_prev_row_count <= 0;
      matmul_11_prev_bat_count <= 0;
      matmul_11_prev_och_count <= 0;
      matmul_11_prev_row_select <= 0;
      matmul_11_out_col_count <= 0;
      matmul_11_out_row_count <= 0;
      matmul_11_out_ram_select <= 0;
      matmul_11_skip_read_filter <= 0;
      matmul_11_skip_read_act <= 0;
      matmul_11_skip_comp <= 0;
      matmul_11_skip_write_out <= 1;
    end else begin
      case(control_matmul_11)
        control_matmul_11_init: begin
          if(main_fsm == 28) begin
            _control_matmul_11_called <= 1;
          end 
          if(main_fsm == 38) begin
            _control_matmul_11_called <= 1;
          end 
          if(main_fsm == 28) begin
            control_matmul_11 <= control_matmul_11_1;
          end 
          if(main_fsm == 38) begin
            control_matmul_11 <= control_matmul_11_1;
          end 
        end
        control_matmul_11_1: begin
          control_matmul_11 <= control_matmul_11_2;
        end
        control_matmul_11_2: begin
          matmul_11_filter_base_offset <= 0;
          matmul_11_filter_page_comp_offset <= 0;
          matmul_11_filter_page_dma_offset <= 0;
          matmul_11_act_base_offset_row <= 0;
          matmul_11_act_base_offset_bat <= 0;
          matmul_11_dma_flag_0 <= 1;
          matmul_11_act_page_comp_offset_0 <= 0;
          matmul_11_act_page_dma_offset_0 <= 0;
          matmul_11_out_base_offset_val <= 0;
          matmul_11_out_base_offset_col <= 0;
          matmul_11_out_base_offset_row <= 0;
          matmul_11_out_base_offset_bat <= 0;
          matmul_11_out_base_offset_och <= 0;
          matmul_11_out_page <= 0;
          matmul_11_out_page_comp_offset <= 0;
          matmul_11_out_page_dma_offset <= 0;
          matmul_11_out_laddr_offset <= 0;
          matmul_11_sync_out_count <= 0;
          matmul_11_write_count <= 0;
          matmul_11_next_out_write_size <= (cparam_matmul_11_max_och_count == 0)? cparam_matmul_11_out_write_size_res : cparam_matmul_11_out_write_size;
          matmul_11_row_count <= 0;
          matmul_11_bat_count <= 0;
          matmul_11_och_count <= 0;
          matmul_11_row_select <= 0;
          matmul_11_prev_row_count <= 0;
          matmul_11_prev_bat_count <= 0;
          matmul_11_prev_och_count <= 0;
          matmul_11_prev_row_select <= 0;
          matmul_11_out_col_count <= 0;
          matmul_11_out_row_count <= 0;
          matmul_11_out_ram_select <= 0;
          matmul_11_skip_read_filter <= 0;
          matmul_11_skip_read_act <= 0;
          matmul_11_skip_comp <= 0;
          matmul_11_skip_write_out <= 1;
          if(_maxi_read_req_idle) begin
            control_matmul_11 <= control_matmul_11_3;
          end 
        end
        control_matmul_11_3: begin
          if(_maxi_read_idle) begin
            control_matmul_11 <= control_matmul_11_4;
          end 
        end
        control_matmul_11_4: begin
          if(_maxi_read_req_idle) begin
            control_matmul_11 <= control_matmul_11_5;
          end 
        end
        control_matmul_11_5: begin
          if(_maxi_read_idle) begin
            control_matmul_11 <= control_matmul_11_6;
          end 
        end
        control_matmul_11_6: begin
          if(cparam_matmul_11_data_stationary == 0) begin
            control_matmul_11 <= control_matmul_11_7;
          end 
          if(cparam_matmul_11_data_stationary == 1) begin
            control_matmul_11 <= control_matmul_11_12;
          end 
        end
        control_matmul_11_7: begin
          control_matmul_11 <= control_matmul_11_8;
          if(matmul_11_skip_read_filter) begin
            control_matmul_11 <= control_matmul_11_11;
          end 
        end
        control_matmul_11_8: begin
          if(_maxi_read_req_idle) begin
            control_matmul_11 <= control_matmul_11_9;
          end 
        end
        control_matmul_11_9: begin
          if(_maxi_read_idle) begin
            control_matmul_11 <= control_matmul_11_10;
          end 
        end
        control_matmul_11_10: begin
          control_matmul_11 <= control_matmul_11_11;
        end
        control_matmul_11_11: begin
          if(cparam_matmul_11_data_stationary == 0) begin
            control_matmul_11 <= control_matmul_11_12;
          end 
          if(cparam_matmul_11_data_stationary == 1) begin
            control_matmul_11 <= control_matmul_11_18;
          end 
        end
        control_matmul_11_12: begin
          control_matmul_11 <= control_matmul_11_13;
          if(matmul_11_skip_read_act) begin
            control_matmul_11 <= control_matmul_11_17;
          end 
        end
        control_matmul_11_13: begin
          control_matmul_11 <= control_matmul_11_14;
          if(matmul_11_mux_dma_pad_mask_0 || !matmul_11_mux_dma_flag_0) begin
            control_matmul_11 <= control_matmul_11_16;
          end 
        end
        control_matmul_11_14: begin
          if(_maxi_read_req_idle) begin
            control_matmul_11 <= control_matmul_11_15;
          end 
        end
        control_matmul_11_15: begin
          if(_maxi_read_idle) begin
            control_matmul_11 <= control_matmul_11_16;
          end 
        end
        control_matmul_11_16: begin
          control_matmul_11 <= control_matmul_11_17;
        end
        control_matmul_11_17: begin
          if(cparam_matmul_11_data_stationary == 0) begin
            control_matmul_11 <= control_matmul_11_18;
          end 
          if(cparam_matmul_11_data_stationary == 1) begin
            control_matmul_11 <= control_matmul_11_7;
          end 
        end
        control_matmul_11_18: begin
          if(_maxi_write_idle) begin
            control_matmul_11 <= control_matmul_11_19;
          end 
        end
        control_matmul_11_19: begin
          if(matmul_11_comp_fsm == 0) begin
            control_matmul_11 <= control_matmul_11_20;
          end 
        end
        control_matmul_11_20: begin
          control_matmul_11 <= control_matmul_11_21;
          if(matmul_11_skip_write_out) begin
            control_matmul_11 <= control_matmul_11_26;
          end 
          if((cparam_matmul_11_data_stationary == 1) && (matmul_11_prev_och_count < cparam_matmul_11_max_och_count)) begin
            control_matmul_11 <= control_matmul_11_26;
          end 
        end
        control_matmul_11_21: begin
          if(matmul_11_sync_comp_count >= matmul_11_sync_out_count + cparam_matmul_11_inc_sync_out) begin
            control_matmul_11 <= control_matmul_11_22;
          end 
        end
        control_matmul_11_22: begin
          if(!matmul_11_dma_out_mask_0) begin
            control_matmul_11 <= control_matmul_11_23;
          end 
          if(matmul_11_dma_out_mask_0) begin
            control_matmul_11 <= control_matmul_11_24;
          end 
        end
        control_matmul_11_23: begin
          if(_maxi_write_req_idle) begin
            control_matmul_11 <= control_matmul_11_24;
          end 
        end
        control_matmul_11_24: begin
          control_matmul_11 <= control_matmul_11_25;
        end
        control_matmul_11_25: begin
          matmul_11_write_count <= matmul_11_write_count + 1;
          if(matmul_11_out_ram_select == 0) begin
            matmul_11_out_laddr_offset <= matmul_11_out_laddr_offset + matmul_11_next_out_write_size;
          end 
          if((cparam_matmul_11_data_stationary == 0) && !cparam_matmul_11_keep_filter) begin
            matmul_11_out_base_offset_col <= matmul_11_out_base_offset_col + cparam_matmul_11_out_col_step;
            matmul_11_out_col_count <= matmul_11_out_col_count + 1;
          end 
          matmul_11_out_ram_select <= matmul_11_out_ram_select + 1;
          if(matmul_11_out_ram_select == 0) begin
            matmul_11_out_ram_select <= 0;
          end 
          matmul_11_sync_out_count <= matmul_11_sync_out_count + cparam_matmul_11_inc_sync_out;
          if((cparam_matmul_11_data_stationary == 0) && !cparam_matmul_11_keep_filter && (matmul_11_write_count >= cparam_matmul_11_out_num_col - 1) || (cparam_matmul_11_data_stationary == 0) && cparam_matmul_11_keep_filter || (cparam_matmul_11_data_stationary == 1)) begin
            matmul_11_sync_out_count <= matmul_11_sync_out_count + (cparam_matmul_11_inc_sync_out + cparam_matmul_11_inc_sync_out_res);
          end 
          if((cparam_matmul_11_data_stationary == 0) && !cparam_matmul_11_keep_filter) begin
            control_matmul_11 <= control_matmul_11_20;
          end 
          if((cparam_matmul_11_data_stationary == 0) && !cparam_matmul_11_keep_filter && (matmul_11_write_count >= cparam_matmul_11_out_num_col - 1) || (cparam_matmul_11_data_stationary == 0) && cparam_matmul_11_keep_filter || (cparam_matmul_11_data_stationary == 1)) begin
            control_matmul_11 <= control_matmul_11_26;
          end 
        end
        control_matmul_11_26: begin
          if(matmul_11_update_filter) begin
            matmul_11_filter_base_offset <= matmul_11_filter_base_offset + cparam_matmul_11_filter_base_step;
          end 
          if((cparam_matmul_11_data_stationary == 1) && (matmul_11_och_count >= cparam_matmul_11_max_och_count)) begin
            matmul_11_filter_base_offset <= 0;
          end 
          if(matmul_11_update_filter) begin
            matmul_11_och_count <= matmul_11_och_count + cparam_matmul_11_och_count_step;
          end 
          if((cparam_matmul_11_data_stationary == 1) && (matmul_11_och_count >= cparam_matmul_11_max_och_count)) begin
            matmul_11_och_count <= 0;
          end 
          if(matmul_11_update_filter) begin
            matmul_11_filter_page_comp_offset <= matmul_11_filter_page_comp_offset + cparam_matmul_11_filter_read_step;
            matmul_11_filter_page_dma_offset <= matmul_11_filter_page_dma_offset + cparam_matmul_11_filter_read_step;
          end 
          if(matmul_11_update_filter && (matmul_11_filter_page_comp_offset + cparam_matmul_11_filter_read_step + cparam_matmul_11_filter_read_step > 32768)) begin
            matmul_11_filter_page_comp_offset <= 0;
            matmul_11_filter_page_dma_offset <= 0;
          end 
          if(matmul_11_update_act) begin
            matmul_11_act_base_offset_row <= matmul_11_act_base_offset_row + cparam_matmul_11_act_row_step;
          end 
          if(matmul_11_update_act && (matmul_11_row_count >= cparam_matmul_11_max_row_count)) begin
            matmul_11_act_base_offset_row <= 0;
            matmul_11_act_base_offset_bat <= matmul_11_act_base_offset_bat + cparam_matmul_11_act_bat_step;
          end 
          if(matmul_11_update_act && (matmul_11_row_count >= cparam_matmul_11_max_row_count) && (matmul_11_bat_count >= cparam_matmul_11_max_bat_count)) begin
            matmul_11_act_base_offset_bat <= 0;
          end 
          if(!matmul_11_update_act) begin
            matmul_11_dma_flag_0 <= 0;
          end 
          if(matmul_11_update_act) begin
            matmul_11_dma_flag_0 <= cparam_matmul_11_dma_flag_conds_0;
          end 
          if(matmul_11_update_act && (matmul_11_row_count >= cparam_matmul_11_max_row_count)) begin
            matmul_11_dma_flag_0 <= 1;
          end 
          if(matmul_11_update_act) begin
            matmul_11_row_count <= matmul_11_row_count + cparam_matmul_11_stride_row_par_row;
          end 
          if(matmul_11_update_act && (matmul_11_row_count >= cparam_matmul_11_max_row_count)) begin
            matmul_11_row_count <= 0;
            matmul_11_bat_count <= matmul_11_bat_count + 1;
          end 
          if(matmul_11_update_act && (matmul_11_row_count >= cparam_matmul_11_max_row_count) && (matmul_11_bat_count >= cparam_matmul_11_max_bat_count)) begin
            matmul_11_bat_count <= 0;
          end 
          if(matmul_11_update_act && (cparam_matmul_11_stride_row_par_row < 1)) begin
            matmul_11_row_select <= matmul_11_row_select + cparam_matmul_11_stride_row_par_row;
            matmul_11_prev_row_select <= matmul_11_row_select;
          end 
          if(matmul_11_update_act && (cparam_matmul_11_stride_row_par_row < 1) && (matmul_11_row_select + cparam_matmul_11_stride_row_par_row >= 1)) begin
            matmul_11_row_select <= matmul_11_row_select - (1 - cparam_matmul_11_stride_row_par_row);
            matmul_11_prev_row_select <= matmul_11_row_select;
          end 
          if(matmul_11_update_act && !(cparam_matmul_11_stride_row_par_row < 1)) begin
            matmul_11_row_select <= 0;
            matmul_11_prev_row_select <= 0;
          end 
          if(matmul_11_update_act && (matmul_11_row_count >= cparam_matmul_11_max_row_count)) begin
            matmul_11_row_select <= 0;
            matmul_11_prev_row_select <= 0;
          end 
          if(matmul_11_update_act && matmul_11_mux_next_dma_flag_0) begin
            matmul_11_act_page_comp_offset_0 <= matmul_11_act_page_comp_offset_0 + cparam_matmul_11_act_read_step;
            matmul_11_act_page_dma_offset_0 <= matmul_11_act_page_dma_offset_0 + cparam_matmul_11_act_read_step;
          end 
          if(matmul_11_update_act && matmul_11_mux_next_dma_flag_0 && (matmul_11_act_page_comp_offset_0 + cparam_matmul_11_act_read_step + cparam_matmul_11_act_read_step > 8192)) begin
            matmul_11_act_page_comp_offset_0 <= 0;
            matmul_11_act_page_dma_offset_0 <= 0;
          end 
          if((cparam_matmul_11_data_stationary == 0) && (matmul_11_row_count >= cparam_matmul_11_max_row_count) && (matmul_11_bat_count >= cparam_matmul_11_max_bat_count) && cparam_matmul_11_keep_input) begin
            matmul_11_act_page_comp_offset_0 <= 0;
            matmul_11_act_page_dma_offset_0 <= 0;
          end 
          matmul_11_next_out_write_size <= (matmul_11_och_count >= cparam_matmul_11_max_och_count)? cparam_matmul_11_out_write_size_res : cparam_matmul_11_out_write_size;
          if(!matmul_11_skip_write_out) begin
            matmul_11_write_count <= 0;
            matmul_11_out_laddr_offset <= 0;
            matmul_11_out_ram_select <= 0;
          end 
          if((cparam_matmul_11_data_stationary == 0) && !matmul_11_skip_write_out) begin
            matmul_11_out_base_offset_col <= 0;
            matmul_11_out_base_offset_row <= matmul_11_out_base_offset_row + cparam_matmul_11_out_row_step;
            matmul_11_out_col_count <= 0;
            matmul_11_out_row_count <= matmul_11_out_row_count + 1;
          end 
          if((cparam_matmul_11_data_stationary == 0) && !matmul_11_skip_write_out && (matmul_11_prev_row_count >= cparam_matmul_11_max_row_count)) begin
            matmul_11_out_base_offset_row <= 0;
            matmul_11_out_base_offset_bat <= matmul_11_out_base_offset_bat + cparam_matmul_11_out_bat_step;
            matmul_11_out_row_count <= 0;
          end 
          if((cparam_matmul_11_data_stationary == 0) && !matmul_11_skip_write_out && (matmul_11_prev_row_count >= cparam_matmul_11_max_row_count) && (matmul_11_prev_bat_count >= cparam_matmul_11_max_bat_count)) begin
            matmul_11_out_base_offset_bat <= 0;
            matmul_11_out_base_offset_och <= matmul_11_out_base_offset_och + cparam_matmul_11_out_och_step;
          end 
          if((cparam_matmul_11_data_stationary == 1) && (matmul_11_prev_och_count >= cparam_matmul_11_max_och_count) && !matmul_11_skip_write_out) begin
            matmul_11_out_base_offset_row <= matmul_11_out_base_offset_row + cparam_matmul_11_out_row_step;
          end 
          if((cparam_matmul_11_data_stationary == 0) && !matmul_11_out_page) begin
            matmul_11_out_page_comp_offset <= 256;
            matmul_11_out_page_dma_offset <= 0;
            matmul_11_out_page <= 1;
          end 
          if((cparam_matmul_11_data_stationary == 0) && matmul_11_out_page) begin
            matmul_11_out_page_comp_offset <= 0;
            matmul_11_out_page_dma_offset <= 256;
            matmul_11_out_page <= 0;
          end 
          if((cparam_matmul_11_data_stationary == 1) && (matmul_11_och_count >= cparam_matmul_11_max_och_count) && !matmul_11_out_page) begin
            matmul_11_out_page_comp_offset <= 256;
            matmul_11_out_page_dma_offset <= 0;
            matmul_11_out_page <= 1;
          end 
          if((cparam_matmul_11_data_stationary == 1) && (matmul_11_och_count >= cparam_matmul_11_max_och_count) && matmul_11_out_page) begin
            matmul_11_out_page_comp_offset <= 0;
            matmul_11_out_page_dma_offset <= 256;
            matmul_11_out_page <= 0;
          end 
          matmul_11_prev_row_count <= matmul_11_row_count;
          matmul_11_prev_bat_count <= matmul_11_bat_count;
          matmul_11_prev_och_count <= matmul_11_och_count;
          if((matmul_11_row_count >= cparam_matmul_11_max_row_count) && (matmul_11_bat_count >= cparam_matmul_11_max_bat_count) && (matmul_11_och_count >= cparam_matmul_11_max_och_count)) begin
            matmul_11_skip_read_filter <= 1;
          end 
          if((cparam_matmul_11_data_stationary == 1) && cparam_matmul_11_keep_filter) begin
            matmul_11_skip_read_filter <= 1;
          end 
          if((matmul_11_row_count >= cparam_matmul_11_max_row_count) && (matmul_11_bat_count >= cparam_matmul_11_max_bat_count) && (matmul_11_och_count >= cparam_matmul_11_max_och_count)) begin
            matmul_11_skip_read_act <= 1;
          end 
          if((cparam_matmul_11_data_stationary == 0) && (matmul_11_row_count >= cparam_matmul_11_max_row_count) && (matmul_11_bat_count >= cparam_matmul_11_max_bat_count) && cparam_matmul_11_keep_input) begin
            matmul_11_skip_read_act <= 1;
          end 
          if((matmul_11_row_count >= cparam_matmul_11_max_row_count) && (matmul_11_bat_count >= cparam_matmul_11_max_bat_count) && (matmul_11_och_count >= cparam_matmul_11_max_och_count)) begin
            matmul_11_skip_comp <= 1;
          end 
          if(matmul_11_skip_write_out && (matmul_11_prev_row_count == 0) && (matmul_11_prev_bat_count == 0) && (matmul_11_prev_och_count == 0)) begin
            matmul_11_skip_write_out <= 0;
          end 
          if(cparam_matmul_11_data_stationary == 0) begin
            control_matmul_11 <= control_matmul_11_12;
          end 
          if((cparam_matmul_11_data_stationary == 0) && (matmul_11_row_count >= cparam_matmul_11_max_row_count) && (matmul_11_bat_count >= cparam_matmul_11_max_bat_count)) begin
            control_matmul_11 <= control_matmul_11_7;
          end 
          if(cparam_matmul_11_data_stationary == 1) begin
            control_matmul_11 <= control_matmul_11_7;
          end 
          if((cparam_matmul_11_data_stationary == 1) && (matmul_11_och_count >= cparam_matmul_11_max_och_count)) begin
            control_matmul_11 <= control_matmul_11_12;
          end 
          if(!matmul_11_skip_write_out && (matmul_11_prev_och_count >= cparam_matmul_11_max_och_count) && (matmul_11_prev_row_count >= cparam_matmul_11_max_row_count) && (matmul_11_prev_bat_count >= cparam_matmul_11_max_bat_count)) begin
            control_matmul_11 <= control_matmul_11_27;
          end 
        end
        control_matmul_11_27: begin
          if(_maxi_write_idle && !_maxi_has_outstanding_write) begin
            control_matmul_11 <= control_matmul_11_28;
          end 
        end
        control_matmul_11_28: begin
          if(main_fsm == 31) begin
            _control_matmul_11_called <= 0;
          end 
          if(main_fsm == 41) begin
            _control_matmul_11_called <= 0;
          end 
          if(main_fsm == 31) begin
            control_matmul_11 <= control_matmul_11_init;
          end 
          if(main_fsm == 41) begin
            control_matmul_11 <= control_matmul_11_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_58_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_58 <= write_burst_packed_fsm_58_init;
      write_burst_packed_addr_1317 <= 0;
      write_burst_packed_stride_1318 <= 0;
      write_burst_packed_length_1319 <= 0;
      write_burst_packed_done_1320 <= 0;
    end else begin
      case(write_burst_packed_fsm_58)
        write_burst_packed_fsm_58_init: begin
          write_burst_packed_addr_1317 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_1318 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_1319 <= _maxi_read_local_size_buf;
          write_burst_packed_done_1320 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 8) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_58 <= write_burst_packed_fsm_58_1;
          end 
        end
        write_burst_packed_fsm_58_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_packed_addr_1317 <= write_burst_packed_addr_1317 + write_burst_packed_stride_1318;
            write_burst_packed_length_1319 <= write_burst_packed_length_1319 - 1;
            write_burst_packed_done_1320 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_packed_length_1319 <= 1)) begin
            write_burst_packed_done_1320 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_packed_done_1320 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_packed_length_1319 <= 1)) begin
            write_burst_packed_fsm_58 <= write_burst_packed_fsm_58_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_packed_fsm_58 <= write_burst_packed_fsm_58_init;
          end 
          if(0) begin
            write_burst_packed_fsm_58 <= write_burst_packed_fsm_58_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_59_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_59 <= write_burst_packed_fsm_59_init;
      write_burst_packed_addr_1330 <= 0;
      write_burst_packed_stride_1331 <= 0;
      write_burst_packed_length_1332 <= 0;
      write_burst_packed_done_1333 <= 0;
    end else begin
      case(write_burst_packed_fsm_59)
        write_burst_packed_fsm_59_init: begin
          write_burst_packed_addr_1330 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_1331 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_1332 <= _maxi_read_local_size_buf;
          write_burst_packed_done_1333 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 9) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_59 <= write_burst_packed_fsm_59_1;
          end 
        end
        write_burst_packed_fsm_59_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_packed_addr_1330 <= write_burst_packed_addr_1330 + write_burst_packed_stride_1331;
            write_burst_packed_length_1332 <= write_burst_packed_length_1332 - 1;
            write_burst_packed_done_1333 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_packed_length_1332 <= 1)) begin
            write_burst_packed_done_1333 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_packed_done_1333 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_packed_length_1332 <= 1)) begin
            write_burst_packed_fsm_59 <= write_burst_packed_fsm_59_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_packed_fsm_59 <= write_burst_packed_fsm_59_init;
          end 
          if(0) begin
            write_burst_packed_fsm_59 <= write_burst_packed_fsm_59_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_60_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_60 <= write_burst_packed_fsm_60_init;
      write_burst_packed_addr_1348 <= 0;
      write_burst_packed_stride_1349 <= 0;
      write_burst_packed_length_1350 <= 0;
      write_burst_packed_done_1351 <= 0;
    end else begin
      case(write_burst_packed_fsm_60)
        write_burst_packed_fsm_60_init: begin
          write_burst_packed_addr_1348 <= _maxi_read_local_addr_buf;
          write_burst_packed_stride_1349 <= _maxi_read_local_stride_buf;
          write_burst_packed_length_1350 <= _maxi_read_local_size_buf;
          write_burst_packed_done_1351 <= 0;
          if((_maxi_read_data_fsm == 1) && (_maxi_read_op_sel_buf == 10) && (_maxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_60 <= write_burst_packed_fsm_60_1;
          end 
        end
        write_burst_packed_fsm_60_1: begin
          if(_maxi_rvalid_sb_0) begin
            write_burst_packed_addr_1348 <= write_burst_packed_addr_1348 + write_burst_packed_stride_1349;
            write_burst_packed_length_1350 <= write_burst_packed_length_1350 - 1;
            write_burst_packed_done_1351 <= 0;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_packed_length_1350 <= 1)) begin
            write_burst_packed_done_1351 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_packed_done_1351 <= 1;
          end 
          if(_maxi_rvalid_sb_0 && (write_burst_packed_length_1350 <= 1)) begin
            write_burst_packed_fsm_60 <= write_burst_packed_fsm_60_init;
          end 
          if(_maxi_rvalid_sb_0 && 0) begin
            write_burst_packed_fsm_60 <= write_burst_packed_fsm_60_init;
          end 
          if(0) begin
            write_burst_packed_fsm_60 <= write_burst_packed_fsm_60_init;
          end 
        end
      endcase
    end
  end

  localparam matmul_11_comp_fsm_1 = 1;
  localparam matmul_11_comp_fsm_2 = 2;
  localparam matmul_11_comp_fsm_3 = 3;
  localparam matmul_11_comp_fsm_4 = 4;
  localparam matmul_11_comp_fsm_5 = 5;
  localparam matmul_11_comp_fsm_6 = 6;

  always @(posedge CLK) begin
    if(RST) begin
      matmul_11_comp_fsm <= matmul_11_comp_fsm_init;
      matmul_11_stream_act_local_0 <= 0;
      matmul_11_stream_out_local_col <= 0;
      matmul_11_stream_out_local_val <= 0;
      matmul_11_col_count <= 0;
      matmul_11_col_select <= 0;
      matmul_11_filter_page_comp_offset_buf <= 0;
      matmul_11_act_page_comp_offset_buf_0 <= 0;
      matmul_11_out_page_comp_offset_buf <= 0;
      matmul_11_row_count_buf <= 0;
      matmul_11_row_select_buf <= 0;
      matmul_11_och_count_buf <= 0;
      matmul_11_next_stream_num_ops <= 0;
      matmul_11_stream_pad_masks <= 0;
      matmul_11_sync_comp_count <= 0;
    end else begin
      if(_stream_matmul_11_sink_stop) begin
        matmul_11_sync_comp_count <= matmul_11_sync_comp_count + 1;
      end 
      if(control_matmul_11 == 6) begin
        matmul_11_sync_comp_count <= 0;
      end 
      case(matmul_11_comp_fsm)
        matmul_11_comp_fsm_init: begin
          if((control_matmul_11 == 19) && !matmul_11_skip_comp) begin
            matmul_11_comp_fsm <= matmul_11_comp_fsm_1;
          end 
        end
        matmul_11_comp_fsm_1: begin
          matmul_11_stream_act_local_0 <= 0;
          if(cparam_matmul_11_stream_act_local_small_flags_0) begin
            matmul_11_stream_act_local_0 <= cparam_matmul_11_stream_act_local_small_offset;
          end 
          if(cparam_matmul_11_stream_act_local_large_flags_0) begin
            matmul_11_stream_act_local_0 <= cparam_matmul_11_stream_act_local_large_offset;
          end 
          matmul_11_stream_out_local_col <= 0;
          if((cparam_matmul_11_data_stationary == 1) && (matmul_11_och_count == 0)) begin
            matmul_11_stream_out_local_val <= 0;
          end 
          matmul_11_col_count <= 0;
          matmul_11_col_select <= cparam_matmul_11_col_select_initval;
          matmul_11_filter_page_comp_offset_buf <= matmul_11_filter_page_comp_offset;
          matmul_11_act_page_comp_offset_buf_0 <= matmul_11_act_page_comp_offset_0;
          matmul_11_out_page_comp_offset_buf <= matmul_11_out_page_comp_offset;
          matmul_11_row_count_buf <= matmul_11_row_count;
          matmul_11_row_select_buf <= matmul_11_row_select;
          matmul_11_och_count_buf <= matmul_11_och_count;
          matmul_11_next_stream_num_ops <= (matmul_11_och_count >= cparam_matmul_11_max_och_count)? cparam_matmul_11_stream_num_ops_res : cparam_matmul_11_stream_num_ops;
          matmul_11_comp_fsm <= matmul_11_comp_fsm_2;
        end
        matmul_11_comp_fsm_2: begin
          matmul_11_stream_pad_masks <= { matmul_11_stream_pad_mask_0_0 };
          matmul_11_comp_fsm <= matmul_11_comp_fsm_3;
        end
        matmul_11_comp_fsm_3: begin
          matmul_11_comp_fsm <= matmul_11_comp_fsm_4;
          matmul_11_comp_fsm <= matmul_11_comp_fsm_4;
          matmul_11_comp_fsm <= matmul_11_comp_fsm_4;
          matmul_11_comp_fsm <= matmul_11_comp_fsm_4;
          matmul_11_comp_fsm <= matmul_11_comp_fsm_4;
          matmul_11_comp_fsm <= matmul_11_comp_fsm_4;
          matmul_11_comp_fsm <= matmul_11_comp_fsm_4;
          matmul_11_comp_fsm <= matmul_11_comp_fsm_4;
          matmul_11_comp_fsm <= matmul_11_comp_fsm_4;
          matmul_11_comp_fsm <= matmul_11_comp_fsm_4;
          matmul_11_comp_fsm <= matmul_11_comp_fsm_4;
          matmul_11_comp_fsm <= matmul_11_comp_fsm_4;
          matmul_11_comp_fsm <= matmul_11_comp_fsm_4;
          matmul_11_comp_fsm <= matmul_11_comp_fsm_4;
          matmul_11_comp_fsm <= matmul_11_comp_fsm_4;
          matmul_11_comp_fsm <= matmul_11_comp_fsm_4;
          matmul_11_comp_fsm <= matmul_11_comp_fsm_4;
          matmul_11_comp_fsm <= matmul_11_comp_fsm_4;
          matmul_11_comp_fsm <= matmul_11_comp_fsm_4;
          matmul_11_comp_fsm <= matmul_11_comp_fsm_4;
          matmul_11_comp_fsm <= matmul_11_comp_fsm_4;
          if(_stream_matmul_11_stream_oready) begin
            matmul_11_comp_fsm <= matmul_11_comp_fsm_4;
          end 
          matmul_11_comp_fsm <= matmul_11_comp_fsm_4;
        end
        matmul_11_comp_fsm_4: begin
          if(!_stream_matmul_11_source_busy) begin
            matmul_11_comp_fsm <= matmul_11_comp_fsm_5;
          end 
        end
        matmul_11_comp_fsm_5: begin
          if(_stream_matmul_11_busy) begin
            matmul_11_comp_fsm <= matmul_11_comp_fsm_6;
          end 
        end
        matmul_11_comp_fsm_6: begin
          if(!((matmul_11_col_select == 0)? cparam_matmul_11_inc_act_laddr_conds_0 : 0)) begin
            matmul_11_stream_act_local_0 <= matmul_11_stream_act_local_0 + cparam_matmul_11_inc_act_laddr_small;
          end 
          if((matmul_11_col_select == 0)? cparam_matmul_11_inc_act_laddr_conds_0 : 0) begin
            matmul_11_stream_act_local_0 <= matmul_11_stream_act_local_0 + cparam_matmul_11_inc_act_laddr_large;
          end 
          if(matmul_11_col_count >= cparam_matmul_11_max_col_count) begin
            matmul_11_stream_act_local_0 <= 0;
          end 
          if((matmul_11_col_count >= cparam_matmul_11_max_col_count) && cparam_matmul_11_stream_act_local_small_flags_0) begin
            matmul_11_stream_act_local_0 <= cparam_matmul_11_stream_act_local_small_offset;
          end 
          if((matmul_11_col_count >= cparam_matmul_11_max_col_count) && cparam_matmul_11_stream_act_local_large_flags_0) begin
            matmul_11_stream_act_local_0 <= cparam_matmul_11_stream_act_local_large_offset;
          end 
          if(cparam_matmul_11_data_stationary == 0) begin
            matmul_11_stream_out_local_col <= matmul_11_stream_out_local_col + matmul_11_next_stream_num_ops;
          end 
          if((cparam_matmul_11_data_stationary == 0) && (matmul_11_col_count >= cparam_matmul_11_max_col_count)) begin
            matmul_11_stream_out_local_col <= 0;
          end 
          if(cparam_matmul_11_data_stationary == 1) begin
            matmul_11_stream_out_local_col <= matmul_11_stream_out_local_col + cparam_matmul_11_inc_out_laddr_col;
          end 
          if((cparam_matmul_11_data_stationary == 1) && (matmul_11_col_count >= cparam_matmul_11_max_col_count)) begin
            matmul_11_stream_out_local_val <= matmul_11_stream_out_local_val + matmul_11_next_stream_num_ops;
            matmul_11_stream_out_local_col <= 0;
          end 
          matmul_11_col_count <= matmul_11_col_count + cparam_matmul_11_stride_col_par_col;
          if(matmul_11_col_count >= cparam_matmul_11_max_col_count) begin
            matmul_11_col_count <= 0;
          end 
          matmul_11_col_select <= matmul_11_col_select + cparam_matmul_11_stride_col_mod_filter_num;
          if(matmul_11_col_select + cparam_matmul_11_stride_col_mod_filter_num >= 1) begin
            matmul_11_col_select <= matmul_11_col_select - cparam_matmul_11_filter_num_col_minus_stride_col_mod;
          end 
          if(matmul_11_col_count >= cparam_matmul_11_max_col_count) begin
            matmul_11_col_select <= cparam_matmul_11_col_select_initval;
          end 
          matmul_11_comp_fsm <= matmul_11_comp_fsm_2;
          if(matmul_11_col_count >= cparam_matmul_11_max_col_count) begin
            matmul_11_comp_fsm <= matmul_11_comp_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_matmul_11_source_7_source_pat_fsm_0_1 = 1;
  localparam _stream_matmul_11_source_7_source_pat_fsm_0_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_matmul_11_source_7_source_pat_fsm_0 <= _stream_matmul_11_source_7_source_pat_fsm_0_init;
    end else begin
      case(_stream_matmul_11_source_7_source_pat_fsm_0)
        _stream_matmul_11_source_7_source_pat_fsm_0_init: begin
          if(_stream_matmul_11_source_start && _stream_matmul_11_source_7_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
            _stream_matmul_11_source_7_source_pat_fsm_0 <= _stream_matmul_11_source_7_source_pat_fsm_0_1;
          end 
        end
        _stream_matmul_11_source_7_source_pat_fsm_0_1: begin
          if(_stream_matmul_11_source_stop && _stream_matmul_11_stream_oready) begin
            _stream_matmul_11_source_7_source_pat_fsm_0 <= _stream_matmul_11_source_7_source_pat_fsm_0_init;
          end 
          if((_source_stream_matmul_11_source_7_pat_count_0 == 0) && (_source_stream_matmul_11_source_7_pat_count_1 == 0) && (_source_stream_matmul_11_source_7_pat_count_2 == 0) && (_source_stream_matmul_11_source_7_pat_count_3 == 0) && _stream_matmul_11_stream_oready) begin
            _stream_matmul_11_source_7_source_pat_fsm_0 <= _stream_matmul_11_source_7_source_pat_fsm_0_2;
          end 
        end
        _stream_matmul_11_source_7_source_pat_fsm_0_2: begin
          if(_stream_matmul_11_stream_oready) begin
            _stream_matmul_11_source_7_source_pat_fsm_0 <= _stream_matmul_11_source_7_source_pat_fsm_0_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_matmul_11_source_9_source_pat_fsm_1_1 = 1;
  localparam _stream_matmul_11_source_9_source_pat_fsm_1_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_matmul_11_source_9_source_pat_fsm_1 <= _stream_matmul_11_source_9_source_pat_fsm_1_init;
    end else begin
      case(_stream_matmul_11_source_9_source_pat_fsm_1)
        _stream_matmul_11_source_9_source_pat_fsm_1_init: begin
          if(_stream_matmul_11_source_start && _stream_matmul_11_source_9_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
            _stream_matmul_11_source_9_source_pat_fsm_1 <= _stream_matmul_11_source_9_source_pat_fsm_1_1;
          end 
        end
        _stream_matmul_11_source_9_source_pat_fsm_1_1: begin
          if(_stream_matmul_11_source_stop && _stream_matmul_11_stream_oready) begin
            _stream_matmul_11_source_9_source_pat_fsm_1 <= _stream_matmul_11_source_9_source_pat_fsm_1_init;
          end 
          if((_source_stream_matmul_11_source_9_pat_count_0 == 0) && (_source_stream_matmul_11_source_9_pat_count_1 == 0) && (_source_stream_matmul_11_source_9_pat_count_2 == 0) && (_source_stream_matmul_11_source_9_pat_count_3 == 0) && _stream_matmul_11_stream_oready) begin
            _stream_matmul_11_source_9_source_pat_fsm_1 <= _stream_matmul_11_source_9_source_pat_fsm_1_2;
          end 
        end
        _stream_matmul_11_source_9_source_pat_fsm_1_2: begin
          if(_stream_matmul_11_stream_oready) begin
            _stream_matmul_11_source_9_source_pat_fsm_1 <= _stream_matmul_11_source_9_source_pat_fsm_1_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_1393 <= 0;
    end else begin
      if(_stream_matmul_11_stream_oready && _stream_matmul_11_source_20_source_ram_renable && (_stream_matmul_11_source_20_source_sel == 3)) begin
        _tmp_1393 <= read_rtl_bank_1392;
      end 
    end
  end

  localparam _stream_matmul_11_source_20_source_pat_fsm_2_1 = 1;
  localparam _stream_matmul_11_source_20_source_pat_fsm_2_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_matmul_11_source_20_source_pat_fsm_2 <= _stream_matmul_11_source_20_source_pat_fsm_2_init;
    end else begin
      case(_stream_matmul_11_source_20_source_pat_fsm_2)
        _stream_matmul_11_source_20_source_pat_fsm_2_init: begin
          if(_stream_matmul_11_source_start && _stream_matmul_11_source_20_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
            _stream_matmul_11_source_20_source_pat_fsm_2 <= _stream_matmul_11_source_20_source_pat_fsm_2_1;
          end 
        end
        _stream_matmul_11_source_20_source_pat_fsm_2_1: begin
          if(_stream_matmul_11_source_stop && _stream_matmul_11_stream_oready) begin
            _stream_matmul_11_source_20_source_pat_fsm_2 <= _stream_matmul_11_source_20_source_pat_fsm_2_init;
          end 
          if((_source_stream_matmul_11_source_20_pat_count_0 == 0) && (_source_stream_matmul_11_source_20_pat_count_1 == 0) && (_source_stream_matmul_11_source_20_pat_count_2 == 0) && (_source_stream_matmul_11_source_20_pat_count_3 == 0) && _stream_matmul_11_stream_oready) begin
            _stream_matmul_11_source_20_source_pat_fsm_2 <= _stream_matmul_11_source_20_source_pat_fsm_2_2;
          end 
        end
        _stream_matmul_11_source_20_source_pat_fsm_2_2: begin
          if(_stream_matmul_11_stream_oready) begin
            _stream_matmul_11_source_20_source_pat_fsm_2 <= _stream_matmul_11_source_20_source_pat_fsm_2_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_matmul_11_source_21_source_pat_fsm_3_1 = 1;
  localparam _stream_matmul_11_source_21_source_pat_fsm_3_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_matmul_11_source_21_source_pat_fsm_3 <= _stream_matmul_11_source_21_source_pat_fsm_3_init;
    end else begin
      case(_stream_matmul_11_source_21_source_pat_fsm_3)
        _stream_matmul_11_source_21_source_pat_fsm_3_init: begin
          if(_stream_matmul_11_source_start && _stream_matmul_11_source_21_source_mode & 5'b10 && _stream_matmul_11_stream_oready) begin
            _stream_matmul_11_source_21_source_pat_fsm_3 <= _stream_matmul_11_source_21_source_pat_fsm_3_1;
          end 
        end
        _stream_matmul_11_source_21_source_pat_fsm_3_1: begin
          if(_stream_matmul_11_source_stop && _stream_matmul_11_stream_oready) begin
            _stream_matmul_11_source_21_source_pat_fsm_3 <= _stream_matmul_11_source_21_source_pat_fsm_3_init;
          end 
          if((_source_stream_matmul_11_source_21_pat_count_0 == 0) && (_source_stream_matmul_11_source_21_pat_count_1 == 0) && (_source_stream_matmul_11_source_21_pat_count_2 == 0) && (_source_stream_matmul_11_source_21_pat_count_3 == 0) && _stream_matmul_11_stream_oready) begin
            _stream_matmul_11_source_21_source_pat_fsm_3 <= _stream_matmul_11_source_21_source_pat_fsm_3_2;
          end 
        end
        _stream_matmul_11_source_21_source_pat_fsm_3_2: begin
          if(_stream_matmul_11_stream_oready) begin
            _stream_matmul_11_source_21_source_pat_fsm_3 <= _stream_matmul_11_source_21_source_pat_fsm_3_init;
          end 
        end
      endcase
    end
  end

  localparam _stream_matmul_11_sink_26_sink_fsm_4_1 = 1;
  localparam _stream_matmul_11_sink_26_sink_fsm_4_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _stream_matmul_11_sink_26_sink_fsm_4 <= _stream_matmul_11_sink_26_sink_fsm_4_init;
    end else begin
      case(_stream_matmul_11_sink_26_sink_fsm_4)
        _stream_matmul_11_sink_26_sink_fsm_4_init: begin
          if(_stream_matmul_11_sink_start && _stream_matmul_11_sink_26_sink_mode & 5'b1 && _stream_matmul_11_stream_oready) begin
            _stream_matmul_11_sink_26_sink_fsm_4 <= _stream_matmul_11_sink_26_sink_fsm_4_1;
          end 
        end
        _stream_matmul_11_sink_26_sink_fsm_4_1: begin
          if(_stream_matmul_11_stream_oready) begin
            _stream_matmul_11_sink_26_sink_fsm_4 <= _stream_matmul_11_sink_26_sink_fsm_4_2;
          end 
        end
        _stream_matmul_11_sink_26_sink_fsm_4_2: begin
          if(stream_matmul_11_sink_27_data && (_stream_matmul_11_sink_26_sink_count == 1) && _stream_matmul_11_stream_oready) begin
            _stream_matmul_11_sink_26_sink_fsm_4 <= _stream_matmul_11_sink_26_sink_fsm_4_init;
          end 
          if(_stream_matmul_11_sink_stop && _stream_matmul_11_stream_oready) begin
            _stream_matmul_11_sink_26_sink_fsm_4 <= _stream_matmul_11_sink_26_sink_fsm_4_init;
          end 
        end
      endcase
    end
  end

  localparam read_burst_packed_fsm_61_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      read_burst_packed_fsm_61 <= read_burst_packed_fsm_61_init;
      read_burst_packed_addr_1632 <= 0;
      read_burst_packed_stride_1633 <= 0;
      read_burst_packed_length_1634 <= 0;
      read_burst_packed_rvalid_1635 <= 0;
      read_burst_packed_rlast_1636 <= 0;
    end else begin
      case(read_burst_packed_fsm_61)
        read_burst_packed_fsm_61_init: begin
          read_burst_packed_addr_1632 <= _maxi_write_local_addr_buf;
          read_burst_packed_stride_1633 <= _maxi_write_local_stride_buf;
          read_burst_packed_length_1634 <= _maxi_write_size_buf;
          read_burst_packed_rvalid_1635 <= 0;
          read_burst_packed_rlast_1636 <= 0;
          if((_maxi_write_data_fsm == 1) && (_maxi_write_op_sel_buf == 3) && (_maxi_write_size_buf > 0)) begin
            read_burst_packed_fsm_61 <= read_burst_packed_fsm_61_1;
          end 
        end
        read_burst_packed_fsm_61_1: begin
          if((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0) && (read_burst_packed_length_1634 > 0)) begin
            read_burst_packed_addr_1632 <= read_burst_packed_addr_1632 + read_burst_packed_stride_1633;
            read_burst_packed_length_1634 <= read_burst_packed_length_1634 - 1;
            read_burst_packed_rvalid_1635 <= 1;
          end 
          if((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0) && (read_burst_packed_length_1634 <= 1)) begin
            read_burst_packed_rlast_1636 <= 1;
          end 
          if(read_burst_packed_rlast_1636 && read_burst_packed_rvalid_1635 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) begin
            read_burst_packed_rvalid_1635 <= 0;
            read_burst_packed_rlast_1636 <= 0;
          end 
          if(0) begin
            read_burst_packed_rvalid_1635 <= 0;
            read_burst_packed_rlast_1636 <= 0;
          end 
          if(read_burst_packed_rlast_1636 && read_burst_packed_rvalid_1635 && ((_maxi_wready_sb_0 || !_maxi_wvalid_sb_0) && (_maxi_write_size_buf > 0))) begin
            read_burst_packed_fsm_61 <= read_burst_packed_fsm_61_init;
          end 
          if(0) begin
            read_burst_packed_fsm_61 <= read_burst_packed_fsm_61_init;
          end 
        end
      endcase
    end
  end


endmodule



module _maxi_read_req_fifo
(
  input CLK,
  input RST,
  input _maxi_read_req_fifo_enq,
  input [137-1:0] _maxi_read_req_fifo_wdata,
  output _maxi_read_req_fifo_full,
  output _maxi_read_req_fifo_almost_full,
  input _maxi_read_req_fifo_deq,
  output [137-1:0] _maxi_read_req_fifo_rdata,
  output _maxi_read_req_fifo_empty,
  output _maxi_read_req_fifo_almost_empty
);

  reg [137-1:0] mem [0:8-1];
  reg [3-1:0] head;
  reg [3-1:0] tail;
  wire is_empty;
  wire is_almost_empty;
  wire is_full;
  wire is_almost_full;
  assign is_empty = head == tail;
  assign is_almost_empty = head == (tail + 1 & 7);
  assign is_full = (head + 1 & 7) == tail;
  assign is_almost_full = (head + 2 & 7) == tail;
  wire [137-1:0] rdata;
  assign _maxi_read_req_fifo_full = is_full;
  assign _maxi_read_req_fifo_almost_full = is_almost_full || is_full;
  assign _maxi_read_req_fifo_empty = is_empty;
  assign _maxi_read_req_fifo_almost_empty = is_almost_empty || is_empty;
  assign rdata = mem[tail];
  assign _maxi_read_req_fifo_rdata = rdata;

  always @(posedge CLK) begin
    if(RST) begin
      head <= 0;
      tail <= 0;
    end else begin
      if(_maxi_read_req_fifo_enq && !is_full) begin
        mem[head] <= _maxi_read_req_fifo_wdata;
        head <= head + 1;
      end 
      if(_maxi_read_req_fifo_deq && !is_empty) begin
        tail <= tail + 1;
      end 
    end
  end


endmodule



module _maxi_write_req_fifo
(
  input CLK,
  input RST,
  input _maxi_write_req_fifo_enq,
  input [137-1:0] _maxi_write_req_fifo_wdata,
  output _maxi_write_req_fifo_full,
  output _maxi_write_req_fifo_almost_full,
  input _maxi_write_req_fifo_deq,
  output [137-1:0] _maxi_write_req_fifo_rdata,
  output _maxi_write_req_fifo_empty,
  output _maxi_write_req_fifo_almost_empty
);

  reg [137-1:0] mem [0:8-1];
  reg [3-1:0] head;
  reg [3-1:0] tail;
  wire is_empty;
  wire is_almost_empty;
  wire is_full;
  wire is_almost_full;
  assign is_empty = head == tail;
  assign is_almost_empty = head == (tail + 1 & 7);
  assign is_full = (head + 1 & 7) == tail;
  assign is_almost_full = (head + 2 & 7) == tail;
  wire [137-1:0] rdata;
  assign _maxi_write_req_fifo_full = is_full;
  assign _maxi_write_req_fifo_almost_full = is_almost_full || is_full;
  assign _maxi_write_req_fifo_empty = is_empty;
  assign _maxi_write_req_fifo_almost_empty = is_almost_empty || is_empty;
  assign rdata = mem[tail];
  assign _maxi_write_req_fifo_rdata = rdata;

  always @(posedge CLK) begin
    if(RST) begin
      head <= 0;
      tail <= 0;
    end else begin
      if(_maxi_write_req_fifo_enq && !is_full) begin
        mem[head] <= _maxi_write_req_fifo_wdata;
        head <= head + 1;
      end 
      if(_maxi_write_req_fifo_deq && !is_empty) begin
        tail <= tail + 1;
      end 
    end
  end


endmodule



module ram_w16_l32768_id0_0
(
  input CLK,
  input [14-1:0] ram_w16_l32768_id0_0_0_addr,
  output [16-1:0] ram_w16_l32768_id0_0_0_rdata,
  input [16-1:0] ram_w16_l32768_id0_0_0_wdata,
  input ram_w16_l32768_id0_0_0_wenable,
  input ram_w16_l32768_id0_0_0_enable,
  input [14-1:0] ram_w16_l32768_id0_0_1_addr,
  output [16-1:0] ram_w16_l32768_id0_0_1_rdata,
  input [16-1:0] ram_w16_l32768_id0_0_1_wdata,
  input ram_w16_l32768_id0_0_1_wenable,
  input ram_w16_l32768_id0_0_1_enable
);

  reg [16-1:0] ram_w16_l32768_id0_0_0_rdata_out;
  assign ram_w16_l32768_id0_0_0_rdata = ram_w16_l32768_id0_0_0_rdata_out;
  reg [16-1:0] ram_w16_l32768_id0_0_1_rdata_out;
  assign ram_w16_l32768_id0_0_1_rdata = ram_w16_l32768_id0_0_1_rdata_out;
  reg [16-1:0] mem [0:16384-1];

  always @(posedge CLK) begin
    if(ram_w16_l32768_id0_0_0_enable) begin
      if(ram_w16_l32768_id0_0_0_wenable) begin
        mem[ram_w16_l32768_id0_0_0_addr] <= ram_w16_l32768_id0_0_0_wdata;
        ram_w16_l32768_id0_0_0_rdata_out <= ram_w16_l32768_id0_0_0_wdata;
      end else begin
        ram_w16_l32768_id0_0_0_rdata_out <= mem[ram_w16_l32768_id0_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l32768_id0_0_1_enable) begin
      if(ram_w16_l32768_id0_0_1_wenable) begin
        mem[ram_w16_l32768_id0_0_1_addr] <= ram_w16_l32768_id0_0_1_wdata;
        ram_w16_l32768_id0_0_1_rdata_out <= ram_w16_l32768_id0_0_1_wdata;
      end else begin
        ram_w16_l32768_id0_0_1_rdata_out <= mem[ram_w16_l32768_id0_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l32768_id0_1
(
  input CLK,
  input [14-1:0] ram_w16_l32768_id0_1_0_addr,
  output [16-1:0] ram_w16_l32768_id0_1_0_rdata,
  input [16-1:0] ram_w16_l32768_id0_1_0_wdata,
  input ram_w16_l32768_id0_1_0_wenable,
  input ram_w16_l32768_id0_1_0_enable,
  input [14-1:0] ram_w16_l32768_id0_1_1_addr,
  output [16-1:0] ram_w16_l32768_id0_1_1_rdata,
  input [16-1:0] ram_w16_l32768_id0_1_1_wdata,
  input ram_w16_l32768_id0_1_1_wenable,
  input ram_w16_l32768_id0_1_1_enable
);

  reg [16-1:0] ram_w16_l32768_id0_1_0_rdata_out;
  assign ram_w16_l32768_id0_1_0_rdata = ram_w16_l32768_id0_1_0_rdata_out;
  reg [16-1:0] ram_w16_l32768_id0_1_1_rdata_out;
  assign ram_w16_l32768_id0_1_1_rdata = ram_w16_l32768_id0_1_1_rdata_out;
  reg [16-1:0] mem [0:16384-1];

  always @(posedge CLK) begin
    if(ram_w16_l32768_id0_1_0_enable) begin
      if(ram_w16_l32768_id0_1_0_wenable) begin
        mem[ram_w16_l32768_id0_1_0_addr] <= ram_w16_l32768_id0_1_0_wdata;
        ram_w16_l32768_id0_1_0_rdata_out <= ram_w16_l32768_id0_1_0_wdata;
      end else begin
        ram_w16_l32768_id0_1_0_rdata_out <= mem[ram_w16_l32768_id0_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l32768_id0_1_1_enable) begin
      if(ram_w16_l32768_id0_1_1_wenable) begin
        mem[ram_w16_l32768_id0_1_1_addr] <= ram_w16_l32768_id0_1_1_wdata;
        ram_w16_l32768_id0_1_1_rdata_out <= ram_w16_l32768_id0_1_1_wdata;
      end else begin
        ram_w16_l32768_id0_1_1_rdata_out <= mem[ram_w16_l32768_id0_1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l8192_id0_0
(
  input CLK,
  input [12-1:0] ram_w16_l8192_id0_0_0_addr,
  output [16-1:0] ram_w16_l8192_id0_0_0_rdata,
  input [16-1:0] ram_w16_l8192_id0_0_0_wdata,
  input ram_w16_l8192_id0_0_0_wenable,
  input ram_w16_l8192_id0_0_0_enable,
  input [12-1:0] ram_w16_l8192_id0_0_1_addr,
  output [16-1:0] ram_w16_l8192_id0_0_1_rdata,
  input [16-1:0] ram_w16_l8192_id0_0_1_wdata,
  input ram_w16_l8192_id0_0_1_wenable,
  input ram_w16_l8192_id0_0_1_enable
);

  reg [16-1:0] ram_w16_l8192_id0_0_0_rdata_out;
  assign ram_w16_l8192_id0_0_0_rdata = ram_w16_l8192_id0_0_0_rdata_out;
  reg [16-1:0] ram_w16_l8192_id0_0_1_rdata_out;
  assign ram_w16_l8192_id0_0_1_rdata = ram_w16_l8192_id0_0_1_rdata_out;
  reg [16-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w16_l8192_id0_0_0_enable) begin
      if(ram_w16_l8192_id0_0_0_wenable) begin
        mem[ram_w16_l8192_id0_0_0_addr] <= ram_w16_l8192_id0_0_0_wdata;
        ram_w16_l8192_id0_0_0_rdata_out <= ram_w16_l8192_id0_0_0_wdata;
      end else begin
        ram_w16_l8192_id0_0_0_rdata_out <= mem[ram_w16_l8192_id0_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l8192_id0_0_1_enable) begin
      if(ram_w16_l8192_id0_0_1_wenable) begin
        mem[ram_w16_l8192_id0_0_1_addr] <= ram_w16_l8192_id0_0_1_wdata;
        ram_w16_l8192_id0_0_1_rdata_out <= ram_w16_l8192_id0_0_1_wdata;
      end else begin
        ram_w16_l8192_id0_0_1_rdata_out <= mem[ram_w16_l8192_id0_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l8192_id0_1
(
  input CLK,
  input [12-1:0] ram_w16_l8192_id0_1_0_addr,
  output [16-1:0] ram_w16_l8192_id0_1_0_rdata,
  input [16-1:0] ram_w16_l8192_id0_1_0_wdata,
  input ram_w16_l8192_id0_1_0_wenable,
  input ram_w16_l8192_id0_1_0_enable,
  input [12-1:0] ram_w16_l8192_id0_1_1_addr,
  output [16-1:0] ram_w16_l8192_id0_1_1_rdata,
  input [16-1:0] ram_w16_l8192_id0_1_1_wdata,
  input ram_w16_l8192_id0_1_1_wenable,
  input ram_w16_l8192_id0_1_1_enable
);

  reg [16-1:0] ram_w16_l8192_id0_1_0_rdata_out;
  assign ram_w16_l8192_id0_1_0_rdata = ram_w16_l8192_id0_1_0_rdata_out;
  reg [16-1:0] ram_w16_l8192_id0_1_1_rdata_out;
  assign ram_w16_l8192_id0_1_1_rdata = ram_w16_l8192_id0_1_1_rdata_out;
  reg [16-1:0] mem [0:4096-1];

  always @(posedge CLK) begin
    if(ram_w16_l8192_id0_1_0_enable) begin
      if(ram_w16_l8192_id0_1_0_wenable) begin
        mem[ram_w16_l8192_id0_1_0_addr] <= ram_w16_l8192_id0_1_0_wdata;
        ram_w16_l8192_id0_1_0_rdata_out <= ram_w16_l8192_id0_1_0_wdata;
      end else begin
        ram_w16_l8192_id0_1_0_rdata_out <= mem[ram_w16_l8192_id0_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l8192_id0_1_1_enable) begin
      if(ram_w16_l8192_id0_1_1_wenable) begin
        mem[ram_w16_l8192_id0_1_1_addr] <= ram_w16_l8192_id0_1_1_wdata;
        ram_w16_l8192_id0_1_1_rdata_out <= ram_w16_l8192_id0_1_1_wdata;
      end else begin
        ram_w16_l8192_id0_1_1_rdata_out <= mem[ram_w16_l8192_id0_1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id0_0
(
  input CLK,
  input [8-1:0] ram_w16_l512_id0_0_0_addr,
  output [16-1:0] ram_w16_l512_id0_0_0_rdata,
  input [16-1:0] ram_w16_l512_id0_0_0_wdata,
  input ram_w16_l512_id0_0_0_wenable,
  input ram_w16_l512_id0_0_0_enable,
  input [8-1:0] ram_w16_l512_id0_0_1_addr,
  output [16-1:0] ram_w16_l512_id0_0_1_rdata,
  input [16-1:0] ram_w16_l512_id0_0_1_wdata,
  input ram_w16_l512_id0_0_1_wenable,
  input ram_w16_l512_id0_0_1_enable
);

  reg [16-1:0] ram_w16_l512_id0_0_0_rdata_out;
  assign ram_w16_l512_id0_0_0_rdata = ram_w16_l512_id0_0_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id0_0_1_rdata_out;
  assign ram_w16_l512_id0_0_1_rdata = ram_w16_l512_id0_0_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id0_0_0_enable) begin
      if(ram_w16_l512_id0_0_0_wenable) begin
        mem[ram_w16_l512_id0_0_0_addr] <= ram_w16_l512_id0_0_0_wdata;
        ram_w16_l512_id0_0_0_rdata_out <= ram_w16_l512_id0_0_0_wdata;
      end else begin
        ram_w16_l512_id0_0_0_rdata_out <= mem[ram_w16_l512_id0_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id0_0_1_enable) begin
      if(ram_w16_l512_id0_0_1_wenable) begin
        mem[ram_w16_l512_id0_0_1_addr] <= ram_w16_l512_id0_0_1_wdata;
        ram_w16_l512_id0_0_1_rdata_out <= ram_w16_l512_id0_0_1_wdata;
      end else begin
        ram_w16_l512_id0_0_1_rdata_out <= mem[ram_w16_l512_id0_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id0_1
(
  input CLK,
  input [8-1:0] ram_w16_l512_id0_1_0_addr,
  output [16-1:0] ram_w16_l512_id0_1_0_rdata,
  input [16-1:0] ram_w16_l512_id0_1_0_wdata,
  input ram_w16_l512_id0_1_0_wenable,
  input ram_w16_l512_id0_1_0_enable,
  input [8-1:0] ram_w16_l512_id0_1_1_addr,
  output [16-1:0] ram_w16_l512_id0_1_1_rdata,
  input [16-1:0] ram_w16_l512_id0_1_1_wdata,
  input ram_w16_l512_id0_1_1_wenable,
  input ram_w16_l512_id0_1_1_enable
);

  reg [16-1:0] ram_w16_l512_id0_1_0_rdata_out;
  assign ram_w16_l512_id0_1_0_rdata = ram_w16_l512_id0_1_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id0_1_1_rdata_out;
  assign ram_w16_l512_id0_1_1_rdata = ram_w16_l512_id0_1_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id0_1_0_enable) begin
      if(ram_w16_l512_id0_1_0_wenable) begin
        mem[ram_w16_l512_id0_1_0_addr] <= ram_w16_l512_id0_1_0_wdata;
        ram_w16_l512_id0_1_0_rdata_out <= ram_w16_l512_id0_1_0_wdata;
      end else begin
        ram_w16_l512_id0_1_0_rdata_out <= mem[ram_w16_l512_id0_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id0_1_1_enable) begin
      if(ram_w16_l512_id0_1_1_wenable) begin
        mem[ram_w16_l512_id0_1_1_addr] <= ram_w16_l512_id0_1_1_wdata;
        ram_w16_l512_id0_1_1_rdata_out <= ram_w16_l512_id0_1_1_wdata;
      end else begin
        ram_w16_l512_id0_1_1_rdata_out <= mem[ram_w16_l512_id0_1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id1_0
(
  input CLK,
  input [8-1:0] ram_w16_l512_id1_0_0_addr,
  output [16-1:0] ram_w16_l512_id1_0_0_rdata,
  input [16-1:0] ram_w16_l512_id1_0_0_wdata,
  input ram_w16_l512_id1_0_0_wenable,
  input ram_w16_l512_id1_0_0_enable,
  input [8-1:0] ram_w16_l512_id1_0_1_addr,
  output [16-1:0] ram_w16_l512_id1_0_1_rdata,
  input [16-1:0] ram_w16_l512_id1_0_1_wdata,
  input ram_w16_l512_id1_0_1_wenable,
  input ram_w16_l512_id1_0_1_enable
);

  reg [16-1:0] ram_w16_l512_id1_0_0_rdata_out;
  assign ram_w16_l512_id1_0_0_rdata = ram_w16_l512_id1_0_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id1_0_1_rdata_out;
  assign ram_w16_l512_id1_0_1_rdata = ram_w16_l512_id1_0_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id1_0_0_enable) begin
      if(ram_w16_l512_id1_0_0_wenable) begin
        mem[ram_w16_l512_id1_0_0_addr] <= ram_w16_l512_id1_0_0_wdata;
        ram_w16_l512_id1_0_0_rdata_out <= ram_w16_l512_id1_0_0_wdata;
      end else begin
        ram_w16_l512_id1_0_0_rdata_out <= mem[ram_w16_l512_id1_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id1_0_1_enable) begin
      if(ram_w16_l512_id1_0_1_wenable) begin
        mem[ram_w16_l512_id1_0_1_addr] <= ram_w16_l512_id1_0_1_wdata;
        ram_w16_l512_id1_0_1_rdata_out <= ram_w16_l512_id1_0_1_wdata;
      end else begin
        ram_w16_l512_id1_0_1_rdata_out <= mem[ram_w16_l512_id1_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id1_1
(
  input CLK,
  input [8-1:0] ram_w16_l512_id1_1_0_addr,
  output [16-1:0] ram_w16_l512_id1_1_0_rdata,
  input [16-1:0] ram_w16_l512_id1_1_0_wdata,
  input ram_w16_l512_id1_1_0_wenable,
  input ram_w16_l512_id1_1_0_enable,
  input [8-1:0] ram_w16_l512_id1_1_1_addr,
  output [16-1:0] ram_w16_l512_id1_1_1_rdata,
  input [16-1:0] ram_w16_l512_id1_1_1_wdata,
  input ram_w16_l512_id1_1_1_wenable,
  input ram_w16_l512_id1_1_1_enable
);

  reg [16-1:0] ram_w16_l512_id1_1_0_rdata_out;
  assign ram_w16_l512_id1_1_0_rdata = ram_w16_l512_id1_1_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id1_1_1_rdata_out;
  assign ram_w16_l512_id1_1_1_rdata = ram_w16_l512_id1_1_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id1_1_0_enable) begin
      if(ram_w16_l512_id1_1_0_wenable) begin
        mem[ram_w16_l512_id1_1_0_addr] <= ram_w16_l512_id1_1_0_wdata;
        ram_w16_l512_id1_1_0_rdata_out <= ram_w16_l512_id1_1_0_wdata;
      end else begin
        ram_w16_l512_id1_1_0_rdata_out <= mem[ram_w16_l512_id1_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id1_1_1_enable) begin
      if(ram_w16_l512_id1_1_1_wenable) begin
        mem[ram_w16_l512_id1_1_1_addr] <= ram_w16_l512_id1_1_1_wdata;
        ram_w16_l512_id1_1_1_rdata_out <= ram_w16_l512_id1_1_1_wdata;
      end else begin
        ram_w16_l512_id1_1_1_rdata_out <= mem[ram_w16_l512_id1_1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id2_0
(
  input CLK,
  input [8-1:0] ram_w16_l512_id2_0_0_addr,
  output [16-1:0] ram_w16_l512_id2_0_0_rdata,
  input [16-1:0] ram_w16_l512_id2_0_0_wdata,
  input ram_w16_l512_id2_0_0_wenable,
  input ram_w16_l512_id2_0_0_enable,
  input [8-1:0] ram_w16_l512_id2_0_1_addr,
  output [16-1:0] ram_w16_l512_id2_0_1_rdata,
  input [16-1:0] ram_w16_l512_id2_0_1_wdata,
  input ram_w16_l512_id2_0_1_wenable,
  input ram_w16_l512_id2_0_1_enable
);

  reg [16-1:0] ram_w16_l512_id2_0_0_rdata_out;
  assign ram_w16_l512_id2_0_0_rdata = ram_w16_l512_id2_0_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id2_0_1_rdata_out;
  assign ram_w16_l512_id2_0_1_rdata = ram_w16_l512_id2_0_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id2_0_0_enable) begin
      if(ram_w16_l512_id2_0_0_wenable) begin
        mem[ram_w16_l512_id2_0_0_addr] <= ram_w16_l512_id2_0_0_wdata;
        ram_w16_l512_id2_0_0_rdata_out <= ram_w16_l512_id2_0_0_wdata;
      end else begin
        ram_w16_l512_id2_0_0_rdata_out <= mem[ram_w16_l512_id2_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id2_0_1_enable) begin
      if(ram_w16_l512_id2_0_1_wenable) begin
        mem[ram_w16_l512_id2_0_1_addr] <= ram_w16_l512_id2_0_1_wdata;
        ram_w16_l512_id2_0_1_rdata_out <= ram_w16_l512_id2_0_1_wdata;
      end else begin
        ram_w16_l512_id2_0_1_rdata_out <= mem[ram_w16_l512_id2_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id2_1
(
  input CLK,
  input [8-1:0] ram_w16_l512_id2_1_0_addr,
  output [16-1:0] ram_w16_l512_id2_1_0_rdata,
  input [16-1:0] ram_w16_l512_id2_1_0_wdata,
  input ram_w16_l512_id2_1_0_wenable,
  input ram_w16_l512_id2_1_0_enable,
  input [8-1:0] ram_w16_l512_id2_1_1_addr,
  output [16-1:0] ram_w16_l512_id2_1_1_rdata,
  input [16-1:0] ram_w16_l512_id2_1_1_wdata,
  input ram_w16_l512_id2_1_1_wenable,
  input ram_w16_l512_id2_1_1_enable
);

  reg [16-1:0] ram_w16_l512_id2_1_0_rdata_out;
  assign ram_w16_l512_id2_1_0_rdata = ram_w16_l512_id2_1_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id2_1_1_rdata_out;
  assign ram_w16_l512_id2_1_1_rdata = ram_w16_l512_id2_1_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id2_1_0_enable) begin
      if(ram_w16_l512_id2_1_0_wenable) begin
        mem[ram_w16_l512_id2_1_0_addr] <= ram_w16_l512_id2_1_0_wdata;
        ram_w16_l512_id2_1_0_rdata_out <= ram_w16_l512_id2_1_0_wdata;
      end else begin
        ram_w16_l512_id2_1_0_rdata_out <= mem[ram_w16_l512_id2_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id2_1_1_enable) begin
      if(ram_w16_l512_id2_1_1_wenable) begin
        mem[ram_w16_l512_id2_1_1_addr] <= ram_w16_l512_id2_1_1_wdata;
        ram_w16_l512_id2_1_1_rdata_out <= ram_w16_l512_id2_1_1_wdata;
      end else begin
        ram_w16_l512_id2_1_1_rdata_out <= mem[ram_w16_l512_id2_1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id3_0
(
  input CLK,
  input [8-1:0] ram_w16_l512_id3_0_0_addr,
  output [16-1:0] ram_w16_l512_id3_0_0_rdata,
  input [16-1:0] ram_w16_l512_id3_0_0_wdata,
  input ram_w16_l512_id3_0_0_wenable,
  input ram_w16_l512_id3_0_0_enable,
  input [8-1:0] ram_w16_l512_id3_0_1_addr,
  output [16-1:0] ram_w16_l512_id3_0_1_rdata,
  input [16-1:0] ram_w16_l512_id3_0_1_wdata,
  input ram_w16_l512_id3_0_1_wenable,
  input ram_w16_l512_id3_0_1_enable
);

  reg [16-1:0] ram_w16_l512_id3_0_0_rdata_out;
  assign ram_w16_l512_id3_0_0_rdata = ram_w16_l512_id3_0_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id3_0_1_rdata_out;
  assign ram_w16_l512_id3_0_1_rdata = ram_w16_l512_id3_0_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id3_0_0_enable) begin
      if(ram_w16_l512_id3_0_0_wenable) begin
        mem[ram_w16_l512_id3_0_0_addr] <= ram_w16_l512_id3_0_0_wdata;
        ram_w16_l512_id3_0_0_rdata_out <= ram_w16_l512_id3_0_0_wdata;
      end else begin
        ram_w16_l512_id3_0_0_rdata_out <= mem[ram_w16_l512_id3_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id3_0_1_enable) begin
      if(ram_w16_l512_id3_0_1_wenable) begin
        mem[ram_w16_l512_id3_0_1_addr] <= ram_w16_l512_id3_0_1_wdata;
        ram_w16_l512_id3_0_1_rdata_out <= ram_w16_l512_id3_0_1_wdata;
      end else begin
        ram_w16_l512_id3_0_1_rdata_out <= mem[ram_w16_l512_id3_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id3_1
(
  input CLK,
  input [8-1:0] ram_w16_l512_id3_1_0_addr,
  output [16-1:0] ram_w16_l512_id3_1_0_rdata,
  input [16-1:0] ram_w16_l512_id3_1_0_wdata,
  input ram_w16_l512_id3_1_0_wenable,
  input ram_w16_l512_id3_1_0_enable,
  input [8-1:0] ram_w16_l512_id3_1_1_addr,
  output [16-1:0] ram_w16_l512_id3_1_1_rdata,
  input [16-1:0] ram_w16_l512_id3_1_1_wdata,
  input ram_w16_l512_id3_1_1_wenable,
  input ram_w16_l512_id3_1_1_enable
);

  reg [16-1:0] ram_w16_l512_id3_1_0_rdata_out;
  assign ram_w16_l512_id3_1_0_rdata = ram_w16_l512_id3_1_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id3_1_1_rdata_out;
  assign ram_w16_l512_id3_1_1_rdata = ram_w16_l512_id3_1_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id3_1_0_enable) begin
      if(ram_w16_l512_id3_1_0_wenable) begin
        mem[ram_w16_l512_id3_1_0_addr] <= ram_w16_l512_id3_1_0_wdata;
        ram_w16_l512_id3_1_0_rdata_out <= ram_w16_l512_id3_1_0_wdata;
      end else begin
        ram_w16_l512_id3_1_0_rdata_out <= mem[ram_w16_l512_id3_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id3_1_1_enable) begin
      if(ram_w16_l512_id3_1_1_wenable) begin
        mem[ram_w16_l512_id3_1_1_addr] <= ram_w16_l512_id3_1_1_wdata;
        ram_w16_l512_id3_1_1_rdata_out <= ram_w16_l512_id3_1_1_wdata;
      end else begin
        ram_w16_l512_id3_1_1_rdata_out <= mem[ram_w16_l512_id3_1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id4_0
(
  input CLK,
  input [8-1:0] ram_w16_l512_id4_0_0_addr,
  output [16-1:0] ram_w16_l512_id4_0_0_rdata,
  input [16-1:0] ram_w16_l512_id4_0_0_wdata,
  input ram_w16_l512_id4_0_0_wenable,
  input ram_w16_l512_id4_0_0_enable,
  input [8-1:0] ram_w16_l512_id4_0_1_addr,
  output [16-1:0] ram_w16_l512_id4_0_1_rdata,
  input [16-1:0] ram_w16_l512_id4_0_1_wdata,
  input ram_w16_l512_id4_0_1_wenable,
  input ram_w16_l512_id4_0_1_enable
);

  reg [16-1:0] ram_w16_l512_id4_0_0_rdata_out;
  assign ram_w16_l512_id4_0_0_rdata = ram_w16_l512_id4_0_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id4_0_1_rdata_out;
  assign ram_w16_l512_id4_0_1_rdata = ram_w16_l512_id4_0_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id4_0_0_enable) begin
      if(ram_w16_l512_id4_0_0_wenable) begin
        mem[ram_w16_l512_id4_0_0_addr] <= ram_w16_l512_id4_0_0_wdata;
        ram_w16_l512_id4_0_0_rdata_out <= ram_w16_l512_id4_0_0_wdata;
      end else begin
        ram_w16_l512_id4_0_0_rdata_out <= mem[ram_w16_l512_id4_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id4_0_1_enable) begin
      if(ram_w16_l512_id4_0_1_wenable) begin
        mem[ram_w16_l512_id4_0_1_addr] <= ram_w16_l512_id4_0_1_wdata;
        ram_w16_l512_id4_0_1_rdata_out <= ram_w16_l512_id4_0_1_wdata;
      end else begin
        ram_w16_l512_id4_0_1_rdata_out <= mem[ram_w16_l512_id4_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id4_1
(
  input CLK,
  input [8-1:0] ram_w16_l512_id4_1_0_addr,
  output [16-1:0] ram_w16_l512_id4_1_0_rdata,
  input [16-1:0] ram_w16_l512_id4_1_0_wdata,
  input ram_w16_l512_id4_1_0_wenable,
  input ram_w16_l512_id4_1_0_enable,
  input [8-1:0] ram_w16_l512_id4_1_1_addr,
  output [16-1:0] ram_w16_l512_id4_1_1_rdata,
  input [16-1:0] ram_w16_l512_id4_1_1_wdata,
  input ram_w16_l512_id4_1_1_wenable,
  input ram_w16_l512_id4_1_1_enable
);

  reg [16-1:0] ram_w16_l512_id4_1_0_rdata_out;
  assign ram_w16_l512_id4_1_0_rdata = ram_w16_l512_id4_1_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id4_1_1_rdata_out;
  assign ram_w16_l512_id4_1_1_rdata = ram_w16_l512_id4_1_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id4_1_0_enable) begin
      if(ram_w16_l512_id4_1_0_wenable) begin
        mem[ram_w16_l512_id4_1_0_addr] <= ram_w16_l512_id4_1_0_wdata;
        ram_w16_l512_id4_1_0_rdata_out <= ram_w16_l512_id4_1_0_wdata;
      end else begin
        ram_w16_l512_id4_1_0_rdata_out <= mem[ram_w16_l512_id4_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id4_1_1_enable) begin
      if(ram_w16_l512_id4_1_1_wenable) begin
        mem[ram_w16_l512_id4_1_1_addr] <= ram_w16_l512_id4_1_1_wdata;
        ram_w16_l512_id4_1_1_rdata_out <= ram_w16_l512_id4_1_1_wdata;
      end else begin
        ram_w16_l512_id4_1_1_rdata_out <= mem[ram_w16_l512_id4_1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id5_0
(
  input CLK,
  input [8-1:0] ram_w16_l512_id5_0_0_addr,
  output [16-1:0] ram_w16_l512_id5_0_0_rdata,
  input [16-1:0] ram_w16_l512_id5_0_0_wdata,
  input ram_w16_l512_id5_0_0_wenable,
  input ram_w16_l512_id5_0_0_enable,
  input [8-1:0] ram_w16_l512_id5_0_1_addr,
  output [16-1:0] ram_w16_l512_id5_0_1_rdata,
  input [16-1:0] ram_w16_l512_id5_0_1_wdata,
  input ram_w16_l512_id5_0_1_wenable,
  input ram_w16_l512_id5_0_1_enable
);

  reg [16-1:0] ram_w16_l512_id5_0_0_rdata_out;
  assign ram_w16_l512_id5_0_0_rdata = ram_w16_l512_id5_0_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id5_0_1_rdata_out;
  assign ram_w16_l512_id5_0_1_rdata = ram_w16_l512_id5_0_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id5_0_0_enable) begin
      if(ram_w16_l512_id5_0_0_wenable) begin
        mem[ram_w16_l512_id5_0_0_addr] <= ram_w16_l512_id5_0_0_wdata;
        ram_w16_l512_id5_0_0_rdata_out <= ram_w16_l512_id5_0_0_wdata;
      end else begin
        ram_w16_l512_id5_0_0_rdata_out <= mem[ram_w16_l512_id5_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id5_0_1_enable) begin
      if(ram_w16_l512_id5_0_1_wenable) begin
        mem[ram_w16_l512_id5_0_1_addr] <= ram_w16_l512_id5_0_1_wdata;
        ram_w16_l512_id5_0_1_rdata_out <= ram_w16_l512_id5_0_1_wdata;
      end else begin
        ram_w16_l512_id5_0_1_rdata_out <= mem[ram_w16_l512_id5_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id5_1
(
  input CLK,
  input [8-1:0] ram_w16_l512_id5_1_0_addr,
  output [16-1:0] ram_w16_l512_id5_1_0_rdata,
  input [16-1:0] ram_w16_l512_id5_1_0_wdata,
  input ram_w16_l512_id5_1_0_wenable,
  input ram_w16_l512_id5_1_0_enable,
  input [8-1:0] ram_w16_l512_id5_1_1_addr,
  output [16-1:0] ram_w16_l512_id5_1_1_rdata,
  input [16-1:0] ram_w16_l512_id5_1_1_wdata,
  input ram_w16_l512_id5_1_1_wenable,
  input ram_w16_l512_id5_1_1_enable
);

  reg [16-1:0] ram_w16_l512_id5_1_0_rdata_out;
  assign ram_w16_l512_id5_1_0_rdata = ram_w16_l512_id5_1_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id5_1_1_rdata_out;
  assign ram_w16_l512_id5_1_1_rdata = ram_w16_l512_id5_1_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id5_1_0_enable) begin
      if(ram_w16_l512_id5_1_0_wenable) begin
        mem[ram_w16_l512_id5_1_0_addr] <= ram_w16_l512_id5_1_0_wdata;
        ram_w16_l512_id5_1_0_rdata_out <= ram_w16_l512_id5_1_0_wdata;
      end else begin
        ram_w16_l512_id5_1_0_rdata_out <= mem[ram_w16_l512_id5_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id5_1_1_enable) begin
      if(ram_w16_l512_id5_1_1_wenable) begin
        mem[ram_w16_l512_id5_1_1_addr] <= ram_w16_l512_id5_1_1_wdata;
        ram_w16_l512_id5_1_1_rdata_out <= ram_w16_l512_id5_1_1_wdata;
      end else begin
        ram_w16_l512_id5_1_1_rdata_out <= mem[ram_w16_l512_id5_1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id6_0
(
  input CLK,
  input [8-1:0] ram_w16_l512_id6_0_0_addr,
  output [16-1:0] ram_w16_l512_id6_0_0_rdata,
  input [16-1:0] ram_w16_l512_id6_0_0_wdata,
  input ram_w16_l512_id6_0_0_wenable,
  input ram_w16_l512_id6_0_0_enable,
  input [8-1:0] ram_w16_l512_id6_0_1_addr,
  output [16-1:0] ram_w16_l512_id6_0_1_rdata,
  input [16-1:0] ram_w16_l512_id6_0_1_wdata,
  input ram_w16_l512_id6_0_1_wenable,
  input ram_w16_l512_id6_0_1_enable
);

  reg [16-1:0] ram_w16_l512_id6_0_0_rdata_out;
  assign ram_w16_l512_id6_0_0_rdata = ram_w16_l512_id6_0_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id6_0_1_rdata_out;
  assign ram_w16_l512_id6_0_1_rdata = ram_w16_l512_id6_0_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id6_0_0_enable) begin
      if(ram_w16_l512_id6_0_0_wenable) begin
        mem[ram_w16_l512_id6_0_0_addr] <= ram_w16_l512_id6_0_0_wdata;
        ram_w16_l512_id6_0_0_rdata_out <= ram_w16_l512_id6_0_0_wdata;
      end else begin
        ram_w16_l512_id6_0_0_rdata_out <= mem[ram_w16_l512_id6_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id6_0_1_enable) begin
      if(ram_w16_l512_id6_0_1_wenable) begin
        mem[ram_w16_l512_id6_0_1_addr] <= ram_w16_l512_id6_0_1_wdata;
        ram_w16_l512_id6_0_1_rdata_out <= ram_w16_l512_id6_0_1_wdata;
      end else begin
        ram_w16_l512_id6_0_1_rdata_out <= mem[ram_w16_l512_id6_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id6_1
(
  input CLK,
  input [8-1:0] ram_w16_l512_id6_1_0_addr,
  output [16-1:0] ram_w16_l512_id6_1_0_rdata,
  input [16-1:0] ram_w16_l512_id6_1_0_wdata,
  input ram_w16_l512_id6_1_0_wenable,
  input ram_w16_l512_id6_1_0_enable,
  input [8-1:0] ram_w16_l512_id6_1_1_addr,
  output [16-1:0] ram_w16_l512_id6_1_1_rdata,
  input [16-1:0] ram_w16_l512_id6_1_1_wdata,
  input ram_w16_l512_id6_1_1_wenable,
  input ram_w16_l512_id6_1_1_enable
);

  reg [16-1:0] ram_w16_l512_id6_1_0_rdata_out;
  assign ram_w16_l512_id6_1_0_rdata = ram_w16_l512_id6_1_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id6_1_1_rdata_out;
  assign ram_w16_l512_id6_1_1_rdata = ram_w16_l512_id6_1_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id6_1_0_enable) begin
      if(ram_w16_l512_id6_1_0_wenable) begin
        mem[ram_w16_l512_id6_1_0_addr] <= ram_w16_l512_id6_1_0_wdata;
        ram_w16_l512_id6_1_0_rdata_out <= ram_w16_l512_id6_1_0_wdata;
      end else begin
        ram_w16_l512_id6_1_0_rdata_out <= mem[ram_w16_l512_id6_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id6_1_1_enable) begin
      if(ram_w16_l512_id6_1_1_wenable) begin
        mem[ram_w16_l512_id6_1_1_addr] <= ram_w16_l512_id6_1_1_wdata;
        ram_w16_l512_id6_1_1_rdata_out <= ram_w16_l512_id6_1_1_wdata;
      end else begin
        ram_w16_l512_id6_1_1_rdata_out <= mem[ram_w16_l512_id6_1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id7_0
(
  input CLK,
  input [8-1:0] ram_w16_l512_id7_0_0_addr,
  output [16-1:0] ram_w16_l512_id7_0_0_rdata,
  input [16-1:0] ram_w16_l512_id7_0_0_wdata,
  input ram_w16_l512_id7_0_0_wenable,
  input ram_w16_l512_id7_0_0_enable,
  input [8-1:0] ram_w16_l512_id7_0_1_addr,
  output [16-1:0] ram_w16_l512_id7_0_1_rdata,
  input [16-1:0] ram_w16_l512_id7_0_1_wdata,
  input ram_w16_l512_id7_0_1_wenable,
  input ram_w16_l512_id7_0_1_enable
);

  reg [16-1:0] ram_w16_l512_id7_0_0_rdata_out;
  assign ram_w16_l512_id7_0_0_rdata = ram_w16_l512_id7_0_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id7_0_1_rdata_out;
  assign ram_w16_l512_id7_0_1_rdata = ram_w16_l512_id7_0_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id7_0_0_enable) begin
      if(ram_w16_l512_id7_0_0_wenable) begin
        mem[ram_w16_l512_id7_0_0_addr] <= ram_w16_l512_id7_0_0_wdata;
        ram_w16_l512_id7_0_0_rdata_out <= ram_w16_l512_id7_0_0_wdata;
      end else begin
        ram_w16_l512_id7_0_0_rdata_out <= mem[ram_w16_l512_id7_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id7_0_1_enable) begin
      if(ram_w16_l512_id7_0_1_wenable) begin
        mem[ram_w16_l512_id7_0_1_addr] <= ram_w16_l512_id7_0_1_wdata;
        ram_w16_l512_id7_0_1_rdata_out <= ram_w16_l512_id7_0_1_wdata;
      end else begin
        ram_w16_l512_id7_0_1_rdata_out <= mem[ram_w16_l512_id7_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id7_1
(
  input CLK,
  input [8-1:0] ram_w16_l512_id7_1_0_addr,
  output [16-1:0] ram_w16_l512_id7_1_0_rdata,
  input [16-1:0] ram_w16_l512_id7_1_0_wdata,
  input ram_w16_l512_id7_1_0_wenable,
  input ram_w16_l512_id7_1_0_enable,
  input [8-1:0] ram_w16_l512_id7_1_1_addr,
  output [16-1:0] ram_w16_l512_id7_1_1_rdata,
  input [16-1:0] ram_w16_l512_id7_1_1_wdata,
  input ram_w16_l512_id7_1_1_wenable,
  input ram_w16_l512_id7_1_1_enable
);

  reg [16-1:0] ram_w16_l512_id7_1_0_rdata_out;
  assign ram_w16_l512_id7_1_0_rdata = ram_w16_l512_id7_1_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id7_1_1_rdata_out;
  assign ram_w16_l512_id7_1_1_rdata = ram_w16_l512_id7_1_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id7_1_0_enable) begin
      if(ram_w16_l512_id7_1_0_wenable) begin
        mem[ram_w16_l512_id7_1_0_addr] <= ram_w16_l512_id7_1_0_wdata;
        ram_w16_l512_id7_1_0_rdata_out <= ram_w16_l512_id7_1_0_wdata;
      end else begin
        ram_w16_l512_id7_1_0_rdata_out <= mem[ram_w16_l512_id7_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id7_1_1_enable) begin
      if(ram_w16_l512_id7_1_1_wenable) begin
        mem[ram_w16_l512_id7_1_1_addr] <= ram_w16_l512_id7_1_1_wdata;
        ram_w16_l512_id7_1_1_rdata_out <= ram_w16_l512_id7_1_1_wdata;
      end else begin
        ram_w16_l512_id7_1_1_rdata_out <= mem[ram_w16_l512_id7_1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id8_0
(
  input CLK,
  input [8-1:0] ram_w16_l512_id8_0_0_addr,
  output [16-1:0] ram_w16_l512_id8_0_0_rdata,
  input [16-1:0] ram_w16_l512_id8_0_0_wdata,
  input ram_w16_l512_id8_0_0_wenable,
  input ram_w16_l512_id8_0_0_enable,
  input [8-1:0] ram_w16_l512_id8_0_1_addr,
  output [16-1:0] ram_w16_l512_id8_0_1_rdata,
  input [16-1:0] ram_w16_l512_id8_0_1_wdata,
  input ram_w16_l512_id8_0_1_wenable,
  input ram_w16_l512_id8_0_1_enable
);

  reg [16-1:0] ram_w16_l512_id8_0_0_rdata_out;
  assign ram_w16_l512_id8_0_0_rdata = ram_w16_l512_id8_0_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id8_0_1_rdata_out;
  assign ram_w16_l512_id8_0_1_rdata = ram_w16_l512_id8_0_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id8_0_0_enable) begin
      if(ram_w16_l512_id8_0_0_wenable) begin
        mem[ram_w16_l512_id8_0_0_addr] <= ram_w16_l512_id8_0_0_wdata;
        ram_w16_l512_id8_0_0_rdata_out <= ram_w16_l512_id8_0_0_wdata;
      end else begin
        ram_w16_l512_id8_0_0_rdata_out <= mem[ram_w16_l512_id8_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id8_0_1_enable) begin
      if(ram_w16_l512_id8_0_1_wenable) begin
        mem[ram_w16_l512_id8_0_1_addr] <= ram_w16_l512_id8_0_1_wdata;
        ram_w16_l512_id8_0_1_rdata_out <= ram_w16_l512_id8_0_1_wdata;
      end else begin
        ram_w16_l512_id8_0_1_rdata_out <= mem[ram_w16_l512_id8_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id8_1
(
  input CLK,
  input [8-1:0] ram_w16_l512_id8_1_0_addr,
  output [16-1:0] ram_w16_l512_id8_1_0_rdata,
  input [16-1:0] ram_w16_l512_id8_1_0_wdata,
  input ram_w16_l512_id8_1_0_wenable,
  input ram_w16_l512_id8_1_0_enable,
  input [8-1:0] ram_w16_l512_id8_1_1_addr,
  output [16-1:0] ram_w16_l512_id8_1_1_rdata,
  input [16-1:0] ram_w16_l512_id8_1_1_wdata,
  input ram_w16_l512_id8_1_1_wenable,
  input ram_w16_l512_id8_1_1_enable
);

  reg [16-1:0] ram_w16_l512_id8_1_0_rdata_out;
  assign ram_w16_l512_id8_1_0_rdata = ram_w16_l512_id8_1_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id8_1_1_rdata_out;
  assign ram_w16_l512_id8_1_1_rdata = ram_w16_l512_id8_1_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id8_1_0_enable) begin
      if(ram_w16_l512_id8_1_0_wenable) begin
        mem[ram_w16_l512_id8_1_0_addr] <= ram_w16_l512_id8_1_0_wdata;
        ram_w16_l512_id8_1_0_rdata_out <= ram_w16_l512_id8_1_0_wdata;
      end else begin
        ram_w16_l512_id8_1_0_rdata_out <= mem[ram_w16_l512_id8_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id8_1_1_enable) begin
      if(ram_w16_l512_id8_1_1_wenable) begin
        mem[ram_w16_l512_id8_1_1_addr] <= ram_w16_l512_id8_1_1_wdata;
        ram_w16_l512_id8_1_1_rdata_out <= ram_w16_l512_id8_1_1_wdata;
      end else begin
        ram_w16_l512_id8_1_1_rdata_out <= mem[ram_w16_l512_id8_1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id9_0
(
  input CLK,
  input [8-1:0] ram_w16_l512_id9_0_0_addr,
  output [16-1:0] ram_w16_l512_id9_0_0_rdata,
  input [16-1:0] ram_w16_l512_id9_0_0_wdata,
  input ram_w16_l512_id9_0_0_wenable,
  input ram_w16_l512_id9_0_0_enable,
  input [8-1:0] ram_w16_l512_id9_0_1_addr,
  output [16-1:0] ram_w16_l512_id9_0_1_rdata,
  input [16-1:0] ram_w16_l512_id9_0_1_wdata,
  input ram_w16_l512_id9_0_1_wenable,
  input ram_w16_l512_id9_0_1_enable
);

  reg [16-1:0] ram_w16_l512_id9_0_0_rdata_out;
  assign ram_w16_l512_id9_0_0_rdata = ram_w16_l512_id9_0_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id9_0_1_rdata_out;
  assign ram_w16_l512_id9_0_1_rdata = ram_w16_l512_id9_0_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id9_0_0_enable) begin
      if(ram_w16_l512_id9_0_0_wenable) begin
        mem[ram_w16_l512_id9_0_0_addr] <= ram_w16_l512_id9_0_0_wdata;
        ram_w16_l512_id9_0_0_rdata_out <= ram_w16_l512_id9_0_0_wdata;
      end else begin
        ram_w16_l512_id9_0_0_rdata_out <= mem[ram_w16_l512_id9_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id9_0_1_enable) begin
      if(ram_w16_l512_id9_0_1_wenable) begin
        mem[ram_w16_l512_id9_0_1_addr] <= ram_w16_l512_id9_0_1_wdata;
        ram_w16_l512_id9_0_1_rdata_out <= ram_w16_l512_id9_0_1_wdata;
      end else begin
        ram_w16_l512_id9_0_1_rdata_out <= mem[ram_w16_l512_id9_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id9_1
(
  input CLK,
  input [8-1:0] ram_w16_l512_id9_1_0_addr,
  output [16-1:0] ram_w16_l512_id9_1_0_rdata,
  input [16-1:0] ram_w16_l512_id9_1_0_wdata,
  input ram_w16_l512_id9_1_0_wenable,
  input ram_w16_l512_id9_1_0_enable,
  input [8-1:0] ram_w16_l512_id9_1_1_addr,
  output [16-1:0] ram_w16_l512_id9_1_1_rdata,
  input [16-1:0] ram_w16_l512_id9_1_1_wdata,
  input ram_w16_l512_id9_1_1_wenable,
  input ram_w16_l512_id9_1_1_enable
);

  reg [16-1:0] ram_w16_l512_id9_1_0_rdata_out;
  assign ram_w16_l512_id9_1_0_rdata = ram_w16_l512_id9_1_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id9_1_1_rdata_out;
  assign ram_w16_l512_id9_1_1_rdata = ram_w16_l512_id9_1_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id9_1_0_enable) begin
      if(ram_w16_l512_id9_1_0_wenable) begin
        mem[ram_w16_l512_id9_1_0_addr] <= ram_w16_l512_id9_1_0_wdata;
        ram_w16_l512_id9_1_0_rdata_out <= ram_w16_l512_id9_1_0_wdata;
      end else begin
        ram_w16_l512_id9_1_0_rdata_out <= mem[ram_w16_l512_id9_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id9_1_1_enable) begin
      if(ram_w16_l512_id9_1_1_wenable) begin
        mem[ram_w16_l512_id9_1_1_addr] <= ram_w16_l512_id9_1_1_wdata;
        ram_w16_l512_id9_1_1_rdata_out <= ram_w16_l512_id9_1_1_wdata;
      end else begin
        ram_w16_l512_id9_1_1_rdata_out <= mem[ram_w16_l512_id9_1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id10_0
(
  input CLK,
  input [8-1:0] ram_w16_l512_id10_0_0_addr,
  output [16-1:0] ram_w16_l512_id10_0_0_rdata,
  input [16-1:0] ram_w16_l512_id10_0_0_wdata,
  input ram_w16_l512_id10_0_0_wenable,
  input ram_w16_l512_id10_0_0_enable,
  input [8-1:0] ram_w16_l512_id10_0_1_addr,
  output [16-1:0] ram_w16_l512_id10_0_1_rdata,
  input [16-1:0] ram_w16_l512_id10_0_1_wdata,
  input ram_w16_l512_id10_0_1_wenable,
  input ram_w16_l512_id10_0_1_enable
);

  reg [16-1:0] ram_w16_l512_id10_0_0_rdata_out;
  assign ram_w16_l512_id10_0_0_rdata = ram_w16_l512_id10_0_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id10_0_1_rdata_out;
  assign ram_w16_l512_id10_0_1_rdata = ram_w16_l512_id10_0_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id10_0_0_enable) begin
      if(ram_w16_l512_id10_0_0_wenable) begin
        mem[ram_w16_l512_id10_0_0_addr] <= ram_w16_l512_id10_0_0_wdata;
        ram_w16_l512_id10_0_0_rdata_out <= ram_w16_l512_id10_0_0_wdata;
      end else begin
        ram_w16_l512_id10_0_0_rdata_out <= mem[ram_w16_l512_id10_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id10_0_1_enable) begin
      if(ram_w16_l512_id10_0_1_wenable) begin
        mem[ram_w16_l512_id10_0_1_addr] <= ram_w16_l512_id10_0_1_wdata;
        ram_w16_l512_id10_0_1_rdata_out <= ram_w16_l512_id10_0_1_wdata;
      end else begin
        ram_w16_l512_id10_0_1_rdata_out <= mem[ram_w16_l512_id10_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id10_1
(
  input CLK,
  input [8-1:0] ram_w16_l512_id10_1_0_addr,
  output [16-1:0] ram_w16_l512_id10_1_0_rdata,
  input [16-1:0] ram_w16_l512_id10_1_0_wdata,
  input ram_w16_l512_id10_1_0_wenable,
  input ram_w16_l512_id10_1_0_enable,
  input [8-1:0] ram_w16_l512_id10_1_1_addr,
  output [16-1:0] ram_w16_l512_id10_1_1_rdata,
  input [16-1:0] ram_w16_l512_id10_1_1_wdata,
  input ram_w16_l512_id10_1_1_wenable,
  input ram_w16_l512_id10_1_1_enable
);

  reg [16-1:0] ram_w16_l512_id10_1_0_rdata_out;
  assign ram_w16_l512_id10_1_0_rdata = ram_w16_l512_id10_1_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id10_1_1_rdata_out;
  assign ram_w16_l512_id10_1_1_rdata = ram_w16_l512_id10_1_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id10_1_0_enable) begin
      if(ram_w16_l512_id10_1_0_wenable) begin
        mem[ram_w16_l512_id10_1_0_addr] <= ram_w16_l512_id10_1_0_wdata;
        ram_w16_l512_id10_1_0_rdata_out <= ram_w16_l512_id10_1_0_wdata;
      end else begin
        ram_w16_l512_id10_1_0_rdata_out <= mem[ram_w16_l512_id10_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id10_1_1_enable) begin
      if(ram_w16_l512_id10_1_1_wenable) begin
        mem[ram_w16_l512_id10_1_1_addr] <= ram_w16_l512_id10_1_1_wdata;
        ram_w16_l512_id10_1_1_rdata_out <= ram_w16_l512_id10_1_1_wdata;
      end else begin
        ram_w16_l512_id10_1_1_rdata_out <= mem[ram_w16_l512_id10_1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id11_0
(
  input CLK,
  input [8-1:0] ram_w16_l512_id11_0_0_addr,
  output [16-1:0] ram_w16_l512_id11_0_0_rdata,
  input [16-1:0] ram_w16_l512_id11_0_0_wdata,
  input ram_w16_l512_id11_0_0_wenable,
  input ram_w16_l512_id11_0_0_enable,
  input [8-1:0] ram_w16_l512_id11_0_1_addr,
  output [16-1:0] ram_w16_l512_id11_0_1_rdata,
  input [16-1:0] ram_w16_l512_id11_0_1_wdata,
  input ram_w16_l512_id11_0_1_wenable,
  input ram_w16_l512_id11_0_1_enable
);

  reg [16-1:0] ram_w16_l512_id11_0_0_rdata_out;
  assign ram_w16_l512_id11_0_0_rdata = ram_w16_l512_id11_0_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id11_0_1_rdata_out;
  assign ram_w16_l512_id11_0_1_rdata = ram_w16_l512_id11_0_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id11_0_0_enable) begin
      if(ram_w16_l512_id11_0_0_wenable) begin
        mem[ram_w16_l512_id11_0_0_addr] <= ram_w16_l512_id11_0_0_wdata;
        ram_w16_l512_id11_0_0_rdata_out <= ram_w16_l512_id11_0_0_wdata;
      end else begin
        ram_w16_l512_id11_0_0_rdata_out <= mem[ram_w16_l512_id11_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id11_0_1_enable) begin
      if(ram_w16_l512_id11_0_1_wenable) begin
        mem[ram_w16_l512_id11_0_1_addr] <= ram_w16_l512_id11_0_1_wdata;
        ram_w16_l512_id11_0_1_rdata_out <= ram_w16_l512_id11_0_1_wdata;
      end else begin
        ram_w16_l512_id11_0_1_rdata_out <= mem[ram_w16_l512_id11_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id11_1
(
  input CLK,
  input [8-1:0] ram_w16_l512_id11_1_0_addr,
  output [16-1:0] ram_w16_l512_id11_1_0_rdata,
  input [16-1:0] ram_w16_l512_id11_1_0_wdata,
  input ram_w16_l512_id11_1_0_wenable,
  input ram_w16_l512_id11_1_0_enable,
  input [8-1:0] ram_w16_l512_id11_1_1_addr,
  output [16-1:0] ram_w16_l512_id11_1_1_rdata,
  input [16-1:0] ram_w16_l512_id11_1_1_wdata,
  input ram_w16_l512_id11_1_1_wenable,
  input ram_w16_l512_id11_1_1_enable
);

  reg [16-1:0] ram_w16_l512_id11_1_0_rdata_out;
  assign ram_w16_l512_id11_1_0_rdata = ram_w16_l512_id11_1_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id11_1_1_rdata_out;
  assign ram_w16_l512_id11_1_1_rdata = ram_w16_l512_id11_1_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id11_1_0_enable) begin
      if(ram_w16_l512_id11_1_0_wenable) begin
        mem[ram_w16_l512_id11_1_0_addr] <= ram_w16_l512_id11_1_0_wdata;
        ram_w16_l512_id11_1_0_rdata_out <= ram_w16_l512_id11_1_0_wdata;
      end else begin
        ram_w16_l512_id11_1_0_rdata_out <= mem[ram_w16_l512_id11_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id11_1_1_enable) begin
      if(ram_w16_l512_id11_1_1_wenable) begin
        mem[ram_w16_l512_id11_1_1_addr] <= ram_w16_l512_id11_1_1_wdata;
        ram_w16_l512_id11_1_1_rdata_out <= ram_w16_l512_id11_1_1_wdata;
      end else begin
        ram_w16_l512_id11_1_1_rdata_out <= mem[ram_w16_l512_id11_1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id12_0
(
  input CLK,
  input [8-1:0] ram_w16_l512_id12_0_0_addr,
  output [16-1:0] ram_w16_l512_id12_0_0_rdata,
  input [16-1:0] ram_w16_l512_id12_0_0_wdata,
  input ram_w16_l512_id12_0_0_wenable,
  input ram_w16_l512_id12_0_0_enable,
  input [8-1:0] ram_w16_l512_id12_0_1_addr,
  output [16-1:0] ram_w16_l512_id12_0_1_rdata,
  input [16-1:0] ram_w16_l512_id12_0_1_wdata,
  input ram_w16_l512_id12_0_1_wenable,
  input ram_w16_l512_id12_0_1_enable
);

  reg [16-1:0] ram_w16_l512_id12_0_0_rdata_out;
  assign ram_w16_l512_id12_0_0_rdata = ram_w16_l512_id12_0_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id12_0_1_rdata_out;
  assign ram_w16_l512_id12_0_1_rdata = ram_w16_l512_id12_0_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id12_0_0_enable) begin
      if(ram_w16_l512_id12_0_0_wenable) begin
        mem[ram_w16_l512_id12_0_0_addr] <= ram_w16_l512_id12_0_0_wdata;
        ram_w16_l512_id12_0_0_rdata_out <= ram_w16_l512_id12_0_0_wdata;
      end else begin
        ram_w16_l512_id12_0_0_rdata_out <= mem[ram_w16_l512_id12_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id12_0_1_enable) begin
      if(ram_w16_l512_id12_0_1_wenable) begin
        mem[ram_w16_l512_id12_0_1_addr] <= ram_w16_l512_id12_0_1_wdata;
        ram_w16_l512_id12_0_1_rdata_out <= ram_w16_l512_id12_0_1_wdata;
      end else begin
        ram_w16_l512_id12_0_1_rdata_out <= mem[ram_w16_l512_id12_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id12_1
(
  input CLK,
  input [8-1:0] ram_w16_l512_id12_1_0_addr,
  output [16-1:0] ram_w16_l512_id12_1_0_rdata,
  input [16-1:0] ram_w16_l512_id12_1_0_wdata,
  input ram_w16_l512_id12_1_0_wenable,
  input ram_w16_l512_id12_1_0_enable,
  input [8-1:0] ram_w16_l512_id12_1_1_addr,
  output [16-1:0] ram_w16_l512_id12_1_1_rdata,
  input [16-1:0] ram_w16_l512_id12_1_1_wdata,
  input ram_w16_l512_id12_1_1_wenable,
  input ram_w16_l512_id12_1_1_enable
);

  reg [16-1:0] ram_w16_l512_id12_1_0_rdata_out;
  assign ram_w16_l512_id12_1_0_rdata = ram_w16_l512_id12_1_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id12_1_1_rdata_out;
  assign ram_w16_l512_id12_1_1_rdata = ram_w16_l512_id12_1_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id12_1_0_enable) begin
      if(ram_w16_l512_id12_1_0_wenable) begin
        mem[ram_w16_l512_id12_1_0_addr] <= ram_w16_l512_id12_1_0_wdata;
        ram_w16_l512_id12_1_0_rdata_out <= ram_w16_l512_id12_1_0_wdata;
      end else begin
        ram_w16_l512_id12_1_0_rdata_out <= mem[ram_w16_l512_id12_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id12_1_1_enable) begin
      if(ram_w16_l512_id12_1_1_wenable) begin
        mem[ram_w16_l512_id12_1_1_addr] <= ram_w16_l512_id12_1_1_wdata;
        ram_w16_l512_id12_1_1_rdata_out <= ram_w16_l512_id12_1_1_wdata;
      end else begin
        ram_w16_l512_id12_1_1_rdata_out <= mem[ram_w16_l512_id12_1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id13_0
(
  input CLK,
  input [8-1:0] ram_w16_l512_id13_0_0_addr,
  output [16-1:0] ram_w16_l512_id13_0_0_rdata,
  input [16-1:0] ram_w16_l512_id13_0_0_wdata,
  input ram_w16_l512_id13_0_0_wenable,
  input ram_w16_l512_id13_0_0_enable,
  input [8-1:0] ram_w16_l512_id13_0_1_addr,
  output [16-1:0] ram_w16_l512_id13_0_1_rdata,
  input [16-1:0] ram_w16_l512_id13_0_1_wdata,
  input ram_w16_l512_id13_0_1_wenable,
  input ram_w16_l512_id13_0_1_enable
);

  reg [16-1:0] ram_w16_l512_id13_0_0_rdata_out;
  assign ram_w16_l512_id13_0_0_rdata = ram_w16_l512_id13_0_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id13_0_1_rdata_out;
  assign ram_w16_l512_id13_0_1_rdata = ram_w16_l512_id13_0_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id13_0_0_enable) begin
      if(ram_w16_l512_id13_0_0_wenable) begin
        mem[ram_w16_l512_id13_0_0_addr] <= ram_w16_l512_id13_0_0_wdata;
        ram_w16_l512_id13_0_0_rdata_out <= ram_w16_l512_id13_0_0_wdata;
      end else begin
        ram_w16_l512_id13_0_0_rdata_out <= mem[ram_w16_l512_id13_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id13_0_1_enable) begin
      if(ram_w16_l512_id13_0_1_wenable) begin
        mem[ram_w16_l512_id13_0_1_addr] <= ram_w16_l512_id13_0_1_wdata;
        ram_w16_l512_id13_0_1_rdata_out <= ram_w16_l512_id13_0_1_wdata;
      end else begin
        ram_w16_l512_id13_0_1_rdata_out <= mem[ram_w16_l512_id13_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id13_1
(
  input CLK,
  input [8-1:0] ram_w16_l512_id13_1_0_addr,
  output [16-1:0] ram_w16_l512_id13_1_0_rdata,
  input [16-1:0] ram_w16_l512_id13_1_0_wdata,
  input ram_w16_l512_id13_1_0_wenable,
  input ram_w16_l512_id13_1_0_enable,
  input [8-1:0] ram_w16_l512_id13_1_1_addr,
  output [16-1:0] ram_w16_l512_id13_1_1_rdata,
  input [16-1:0] ram_w16_l512_id13_1_1_wdata,
  input ram_w16_l512_id13_1_1_wenable,
  input ram_w16_l512_id13_1_1_enable
);

  reg [16-1:0] ram_w16_l512_id13_1_0_rdata_out;
  assign ram_w16_l512_id13_1_0_rdata = ram_w16_l512_id13_1_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id13_1_1_rdata_out;
  assign ram_w16_l512_id13_1_1_rdata = ram_w16_l512_id13_1_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id13_1_0_enable) begin
      if(ram_w16_l512_id13_1_0_wenable) begin
        mem[ram_w16_l512_id13_1_0_addr] <= ram_w16_l512_id13_1_0_wdata;
        ram_w16_l512_id13_1_0_rdata_out <= ram_w16_l512_id13_1_0_wdata;
      end else begin
        ram_w16_l512_id13_1_0_rdata_out <= mem[ram_w16_l512_id13_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id13_1_1_enable) begin
      if(ram_w16_l512_id13_1_1_wenable) begin
        mem[ram_w16_l512_id13_1_1_addr] <= ram_w16_l512_id13_1_1_wdata;
        ram_w16_l512_id13_1_1_rdata_out <= ram_w16_l512_id13_1_1_wdata;
      end else begin
        ram_w16_l512_id13_1_1_rdata_out <= mem[ram_w16_l512_id13_1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id14_0
(
  input CLK,
  input [8-1:0] ram_w16_l512_id14_0_0_addr,
  output [16-1:0] ram_w16_l512_id14_0_0_rdata,
  input [16-1:0] ram_w16_l512_id14_0_0_wdata,
  input ram_w16_l512_id14_0_0_wenable,
  input ram_w16_l512_id14_0_0_enable,
  input [8-1:0] ram_w16_l512_id14_0_1_addr,
  output [16-1:0] ram_w16_l512_id14_0_1_rdata,
  input [16-1:0] ram_w16_l512_id14_0_1_wdata,
  input ram_w16_l512_id14_0_1_wenable,
  input ram_w16_l512_id14_0_1_enable
);

  reg [16-1:0] ram_w16_l512_id14_0_0_rdata_out;
  assign ram_w16_l512_id14_0_0_rdata = ram_w16_l512_id14_0_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id14_0_1_rdata_out;
  assign ram_w16_l512_id14_0_1_rdata = ram_w16_l512_id14_0_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id14_0_0_enable) begin
      if(ram_w16_l512_id14_0_0_wenable) begin
        mem[ram_w16_l512_id14_0_0_addr] <= ram_w16_l512_id14_0_0_wdata;
        ram_w16_l512_id14_0_0_rdata_out <= ram_w16_l512_id14_0_0_wdata;
      end else begin
        ram_w16_l512_id14_0_0_rdata_out <= mem[ram_w16_l512_id14_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id14_0_1_enable) begin
      if(ram_w16_l512_id14_0_1_wenable) begin
        mem[ram_w16_l512_id14_0_1_addr] <= ram_w16_l512_id14_0_1_wdata;
        ram_w16_l512_id14_0_1_rdata_out <= ram_w16_l512_id14_0_1_wdata;
      end else begin
        ram_w16_l512_id14_0_1_rdata_out <= mem[ram_w16_l512_id14_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id14_1
(
  input CLK,
  input [8-1:0] ram_w16_l512_id14_1_0_addr,
  output [16-1:0] ram_w16_l512_id14_1_0_rdata,
  input [16-1:0] ram_w16_l512_id14_1_0_wdata,
  input ram_w16_l512_id14_1_0_wenable,
  input ram_w16_l512_id14_1_0_enable,
  input [8-1:0] ram_w16_l512_id14_1_1_addr,
  output [16-1:0] ram_w16_l512_id14_1_1_rdata,
  input [16-1:0] ram_w16_l512_id14_1_1_wdata,
  input ram_w16_l512_id14_1_1_wenable,
  input ram_w16_l512_id14_1_1_enable
);

  reg [16-1:0] ram_w16_l512_id14_1_0_rdata_out;
  assign ram_w16_l512_id14_1_0_rdata = ram_w16_l512_id14_1_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id14_1_1_rdata_out;
  assign ram_w16_l512_id14_1_1_rdata = ram_w16_l512_id14_1_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id14_1_0_enable) begin
      if(ram_w16_l512_id14_1_0_wenable) begin
        mem[ram_w16_l512_id14_1_0_addr] <= ram_w16_l512_id14_1_0_wdata;
        ram_w16_l512_id14_1_0_rdata_out <= ram_w16_l512_id14_1_0_wdata;
      end else begin
        ram_w16_l512_id14_1_0_rdata_out <= mem[ram_w16_l512_id14_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id14_1_1_enable) begin
      if(ram_w16_l512_id14_1_1_wenable) begin
        mem[ram_w16_l512_id14_1_1_addr] <= ram_w16_l512_id14_1_1_wdata;
        ram_w16_l512_id14_1_1_rdata_out <= ram_w16_l512_id14_1_1_wdata;
      end else begin
        ram_w16_l512_id14_1_1_rdata_out <= mem[ram_w16_l512_id14_1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id15_0
(
  input CLK,
  input [8-1:0] ram_w16_l512_id15_0_0_addr,
  output [16-1:0] ram_w16_l512_id15_0_0_rdata,
  input [16-1:0] ram_w16_l512_id15_0_0_wdata,
  input ram_w16_l512_id15_0_0_wenable,
  input ram_w16_l512_id15_0_0_enable,
  input [8-1:0] ram_w16_l512_id15_0_1_addr,
  output [16-1:0] ram_w16_l512_id15_0_1_rdata,
  input [16-1:0] ram_w16_l512_id15_0_1_wdata,
  input ram_w16_l512_id15_0_1_wenable,
  input ram_w16_l512_id15_0_1_enable
);

  reg [16-1:0] ram_w16_l512_id15_0_0_rdata_out;
  assign ram_w16_l512_id15_0_0_rdata = ram_w16_l512_id15_0_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id15_0_1_rdata_out;
  assign ram_w16_l512_id15_0_1_rdata = ram_w16_l512_id15_0_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id15_0_0_enable) begin
      if(ram_w16_l512_id15_0_0_wenable) begin
        mem[ram_w16_l512_id15_0_0_addr] <= ram_w16_l512_id15_0_0_wdata;
        ram_w16_l512_id15_0_0_rdata_out <= ram_w16_l512_id15_0_0_wdata;
      end else begin
        ram_w16_l512_id15_0_0_rdata_out <= mem[ram_w16_l512_id15_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id15_0_1_enable) begin
      if(ram_w16_l512_id15_0_1_wenable) begin
        mem[ram_w16_l512_id15_0_1_addr] <= ram_w16_l512_id15_0_1_wdata;
        ram_w16_l512_id15_0_1_rdata_out <= ram_w16_l512_id15_0_1_wdata;
      end else begin
        ram_w16_l512_id15_0_1_rdata_out <= mem[ram_w16_l512_id15_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id15_1
(
  input CLK,
  input [8-1:0] ram_w16_l512_id15_1_0_addr,
  output [16-1:0] ram_w16_l512_id15_1_0_rdata,
  input [16-1:0] ram_w16_l512_id15_1_0_wdata,
  input ram_w16_l512_id15_1_0_wenable,
  input ram_w16_l512_id15_1_0_enable,
  input [8-1:0] ram_w16_l512_id15_1_1_addr,
  output [16-1:0] ram_w16_l512_id15_1_1_rdata,
  input [16-1:0] ram_w16_l512_id15_1_1_wdata,
  input ram_w16_l512_id15_1_1_wenable,
  input ram_w16_l512_id15_1_1_enable
);

  reg [16-1:0] ram_w16_l512_id15_1_0_rdata_out;
  assign ram_w16_l512_id15_1_0_rdata = ram_w16_l512_id15_1_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id15_1_1_rdata_out;
  assign ram_w16_l512_id15_1_1_rdata = ram_w16_l512_id15_1_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id15_1_0_enable) begin
      if(ram_w16_l512_id15_1_0_wenable) begin
        mem[ram_w16_l512_id15_1_0_addr] <= ram_w16_l512_id15_1_0_wdata;
        ram_w16_l512_id15_1_0_rdata_out <= ram_w16_l512_id15_1_0_wdata;
      end else begin
        ram_w16_l512_id15_1_0_rdata_out <= mem[ram_w16_l512_id15_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id15_1_1_enable) begin
      if(ram_w16_l512_id15_1_1_wenable) begin
        mem[ram_w16_l512_id15_1_1_addr] <= ram_w16_l512_id15_1_1_wdata;
        ram_w16_l512_id15_1_1_rdata_out <= ram_w16_l512_id15_1_1_wdata;
      end else begin
        ram_w16_l512_id15_1_1_rdata_out <= mem[ram_w16_l512_id15_1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id16_0
(
  input CLK,
  input [8-1:0] ram_w16_l512_id16_0_0_addr,
  output [16-1:0] ram_w16_l512_id16_0_0_rdata,
  input [16-1:0] ram_w16_l512_id16_0_0_wdata,
  input ram_w16_l512_id16_0_0_wenable,
  input ram_w16_l512_id16_0_0_enable,
  input [8-1:0] ram_w16_l512_id16_0_1_addr,
  output [16-1:0] ram_w16_l512_id16_0_1_rdata,
  input [16-1:0] ram_w16_l512_id16_0_1_wdata,
  input ram_w16_l512_id16_0_1_wenable,
  input ram_w16_l512_id16_0_1_enable
);

  reg [16-1:0] ram_w16_l512_id16_0_0_rdata_out;
  assign ram_w16_l512_id16_0_0_rdata = ram_w16_l512_id16_0_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id16_0_1_rdata_out;
  assign ram_w16_l512_id16_0_1_rdata = ram_w16_l512_id16_0_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id16_0_0_enable) begin
      if(ram_w16_l512_id16_0_0_wenable) begin
        mem[ram_w16_l512_id16_0_0_addr] <= ram_w16_l512_id16_0_0_wdata;
        ram_w16_l512_id16_0_0_rdata_out <= ram_w16_l512_id16_0_0_wdata;
      end else begin
        ram_w16_l512_id16_0_0_rdata_out <= mem[ram_w16_l512_id16_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id16_0_1_enable) begin
      if(ram_w16_l512_id16_0_1_wenable) begin
        mem[ram_w16_l512_id16_0_1_addr] <= ram_w16_l512_id16_0_1_wdata;
        ram_w16_l512_id16_0_1_rdata_out <= ram_w16_l512_id16_0_1_wdata;
      end else begin
        ram_w16_l512_id16_0_1_rdata_out <= mem[ram_w16_l512_id16_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id16_1
(
  input CLK,
  input [8-1:0] ram_w16_l512_id16_1_0_addr,
  output [16-1:0] ram_w16_l512_id16_1_0_rdata,
  input [16-1:0] ram_w16_l512_id16_1_0_wdata,
  input ram_w16_l512_id16_1_0_wenable,
  input ram_w16_l512_id16_1_0_enable,
  input [8-1:0] ram_w16_l512_id16_1_1_addr,
  output [16-1:0] ram_w16_l512_id16_1_1_rdata,
  input [16-1:0] ram_w16_l512_id16_1_1_wdata,
  input ram_w16_l512_id16_1_1_wenable,
  input ram_w16_l512_id16_1_1_enable
);

  reg [16-1:0] ram_w16_l512_id16_1_0_rdata_out;
  assign ram_w16_l512_id16_1_0_rdata = ram_w16_l512_id16_1_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id16_1_1_rdata_out;
  assign ram_w16_l512_id16_1_1_rdata = ram_w16_l512_id16_1_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id16_1_0_enable) begin
      if(ram_w16_l512_id16_1_0_wenable) begin
        mem[ram_w16_l512_id16_1_0_addr] <= ram_w16_l512_id16_1_0_wdata;
        ram_w16_l512_id16_1_0_rdata_out <= ram_w16_l512_id16_1_0_wdata;
      end else begin
        ram_w16_l512_id16_1_0_rdata_out <= mem[ram_w16_l512_id16_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id16_1_1_enable) begin
      if(ram_w16_l512_id16_1_1_wenable) begin
        mem[ram_w16_l512_id16_1_1_addr] <= ram_w16_l512_id16_1_1_wdata;
        ram_w16_l512_id16_1_1_rdata_out <= ram_w16_l512_id16_1_1_wdata;
      end else begin
        ram_w16_l512_id16_1_1_rdata_out <= mem[ram_w16_l512_id16_1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id17_0
(
  input CLK,
  input [8-1:0] ram_w16_l512_id17_0_0_addr,
  output [16-1:0] ram_w16_l512_id17_0_0_rdata,
  input [16-1:0] ram_w16_l512_id17_0_0_wdata,
  input ram_w16_l512_id17_0_0_wenable,
  input ram_w16_l512_id17_0_0_enable,
  input [8-1:0] ram_w16_l512_id17_0_1_addr,
  output [16-1:0] ram_w16_l512_id17_0_1_rdata,
  input [16-1:0] ram_w16_l512_id17_0_1_wdata,
  input ram_w16_l512_id17_0_1_wenable,
  input ram_w16_l512_id17_0_1_enable
);

  reg [16-1:0] ram_w16_l512_id17_0_0_rdata_out;
  assign ram_w16_l512_id17_0_0_rdata = ram_w16_l512_id17_0_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id17_0_1_rdata_out;
  assign ram_w16_l512_id17_0_1_rdata = ram_w16_l512_id17_0_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id17_0_0_enable) begin
      if(ram_w16_l512_id17_0_0_wenable) begin
        mem[ram_w16_l512_id17_0_0_addr] <= ram_w16_l512_id17_0_0_wdata;
        ram_w16_l512_id17_0_0_rdata_out <= ram_w16_l512_id17_0_0_wdata;
      end else begin
        ram_w16_l512_id17_0_0_rdata_out <= mem[ram_w16_l512_id17_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id17_0_1_enable) begin
      if(ram_w16_l512_id17_0_1_wenable) begin
        mem[ram_w16_l512_id17_0_1_addr] <= ram_w16_l512_id17_0_1_wdata;
        ram_w16_l512_id17_0_1_rdata_out <= ram_w16_l512_id17_0_1_wdata;
      end else begin
        ram_w16_l512_id17_0_1_rdata_out <= mem[ram_w16_l512_id17_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id17_1
(
  input CLK,
  input [8-1:0] ram_w16_l512_id17_1_0_addr,
  output [16-1:0] ram_w16_l512_id17_1_0_rdata,
  input [16-1:0] ram_w16_l512_id17_1_0_wdata,
  input ram_w16_l512_id17_1_0_wenable,
  input ram_w16_l512_id17_1_0_enable,
  input [8-1:0] ram_w16_l512_id17_1_1_addr,
  output [16-1:0] ram_w16_l512_id17_1_1_rdata,
  input [16-1:0] ram_w16_l512_id17_1_1_wdata,
  input ram_w16_l512_id17_1_1_wenable,
  input ram_w16_l512_id17_1_1_enable
);

  reg [16-1:0] ram_w16_l512_id17_1_0_rdata_out;
  assign ram_w16_l512_id17_1_0_rdata = ram_w16_l512_id17_1_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id17_1_1_rdata_out;
  assign ram_w16_l512_id17_1_1_rdata = ram_w16_l512_id17_1_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id17_1_0_enable) begin
      if(ram_w16_l512_id17_1_0_wenable) begin
        mem[ram_w16_l512_id17_1_0_addr] <= ram_w16_l512_id17_1_0_wdata;
        ram_w16_l512_id17_1_0_rdata_out <= ram_w16_l512_id17_1_0_wdata;
      end else begin
        ram_w16_l512_id17_1_0_rdata_out <= mem[ram_w16_l512_id17_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id17_1_1_enable) begin
      if(ram_w16_l512_id17_1_1_wenable) begin
        mem[ram_w16_l512_id17_1_1_addr] <= ram_w16_l512_id17_1_1_wdata;
        ram_w16_l512_id17_1_1_rdata_out <= ram_w16_l512_id17_1_1_wdata;
      end else begin
        ram_w16_l512_id17_1_1_rdata_out <= mem[ram_w16_l512_id17_1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id18_0
(
  input CLK,
  input [8-1:0] ram_w16_l512_id18_0_0_addr,
  output [16-1:0] ram_w16_l512_id18_0_0_rdata,
  input [16-1:0] ram_w16_l512_id18_0_0_wdata,
  input ram_w16_l512_id18_0_0_wenable,
  input ram_w16_l512_id18_0_0_enable,
  input [8-1:0] ram_w16_l512_id18_0_1_addr,
  output [16-1:0] ram_w16_l512_id18_0_1_rdata,
  input [16-1:0] ram_w16_l512_id18_0_1_wdata,
  input ram_w16_l512_id18_0_1_wenable,
  input ram_w16_l512_id18_0_1_enable
);

  reg [16-1:0] ram_w16_l512_id18_0_0_rdata_out;
  assign ram_w16_l512_id18_0_0_rdata = ram_w16_l512_id18_0_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id18_0_1_rdata_out;
  assign ram_w16_l512_id18_0_1_rdata = ram_w16_l512_id18_0_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id18_0_0_enable) begin
      if(ram_w16_l512_id18_0_0_wenable) begin
        mem[ram_w16_l512_id18_0_0_addr] <= ram_w16_l512_id18_0_0_wdata;
        ram_w16_l512_id18_0_0_rdata_out <= ram_w16_l512_id18_0_0_wdata;
      end else begin
        ram_w16_l512_id18_0_0_rdata_out <= mem[ram_w16_l512_id18_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id18_0_1_enable) begin
      if(ram_w16_l512_id18_0_1_wenable) begin
        mem[ram_w16_l512_id18_0_1_addr] <= ram_w16_l512_id18_0_1_wdata;
        ram_w16_l512_id18_0_1_rdata_out <= ram_w16_l512_id18_0_1_wdata;
      end else begin
        ram_w16_l512_id18_0_1_rdata_out <= mem[ram_w16_l512_id18_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id18_1
(
  input CLK,
  input [8-1:0] ram_w16_l512_id18_1_0_addr,
  output [16-1:0] ram_w16_l512_id18_1_0_rdata,
  input [16-1:0] ram_w16_l512_id18_1_0_wdata,
  input ram_w16_l512_id18_1_0_wenable,
  input ram_w16_l512_id18_1_0_enable,
  input [8-1:0] ram_w16_l512_id18_1_1_addr,
  output [16-1:0] ram_w16_l512_id18_1_1_rdata,
  input [16-1:0] ram_w16_l512_id18_1_1_wdata,
  input ram_w16_l512_id18_1_1_wenable,
  input ram_w16_l512_id18_1_1_enable
);

  reg [16-1:0] ram_w16_l512_id18_1_0_rdata_out;
  assign ram_w16_l512_id18_1_0_rdata = ram_w16_l512_id18_1_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id18_1_1_rdata_out;
  assign ram_w16_l512_id18_1_1_rdata = ram_w16_l512_id18_1_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id18_1_0_enable) begin
      if(ram_w16_l512_id18_1_0_wenable) begin
        mem[ram_w16_l512_id18_1_0_addr] <= ram_w16_l512_id18_1_0_wdata;
        ram_w16_l512_id18_1_0_rdata_out <= ram_w16_l512_id18_1_0_wdata;
      end else begin
        ram_w16_l512_id18_1_0_rdata_out <= mem[ram_w16_l512_id18_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id18_1_1_enable) begin
      if(ram_w16_l512_id18_1_1_wenable) begin
        mem[ram_w16_l512_id18_1_1_addr] <= ram_w16_l512_id18_1_1_wdata;
        ram_w16_l512_id18_1_1_rdata_out <= ram_w16_l512_id18_1_1_wdata;
      end else begin
        ram_w16_l512_id18_1_1_rdata_out <= mem[ram_w16_l512_id18_1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id19_0
(
  input CLK,
  input [8-1:0] ram_w16_l512_id19_0_0_addr,
  output [16-1:0] ram_w16_l512_id19_0_0_rdata,
  input [16-1:0] ram_w16_l512_id19_0_0_wdata,
  input ram_w16_l512_id19_0_0_wenable,
  input ram_w16_l512_id19_0_0_enable,
  input [8-1:0] ram_w16_l512_id19_0_1_addr,
  output [16-1:0] ram_w16_l512_id19_0_1_rdata,
  input [16-1:0] ram_w16_l512_id19_0_1_wdata,
  input ram_w16_l512_id19_0_1_wenable,
  input ram_w16_l512_id19_0_1_enable
);

  reg [16-1:0] ram_w16_l512_id19_0_0_rdata_out;
  assign ram_w16_l512_id19_0_0_rdata = ram_w16_l512_id19_0_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id19_0_1_rdata_out;
  assign ram_w16_l512_id19_0_1_rdata = ram_w16_l512_id19_0_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id19_0_0_enable) begin
      if(ram_w16_l512_id19_0_0_wenable) begin
        mem[ram_w16_l512_id19_0_0_addr] <= ram_w16_l512_id19_0_0_wdata;
        ram_w16_l512_id19_0_0_rdata_out <= ram_w16_l512_id19_0_0_wdata;
      end else begin
        ram_w16_l512_id19_0_0_rdata_out <= mem[ram_w16_l512_id19_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id19_0_1_enable) begin
      if(ram_w16_l512_id19_0_1_wenable) begin
        mem[ram_w16_l512_id19_0_1_addr] <= ram_w16_l512_id19_0_1_wdata;
        ram_w16_l512_id19_0_1_rdata_out <= ram_w16_l512_id19_0_1_wdata;
      end else begin
        ram_w16_l512_id19_0_1_rdata_out <= mem[ram_w16_l512_id19_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id19_1
(
  input CLK,
  input [8-1:0] ram_w16_l512_id19_1_0_addr,
  output [16-1:0] ram_w16_l512_id19_1_0_rdata,
  input [16-1:0] ram_w16_l512_id19_1_0_wdata,
  input ram_w16_l512_id19_1_0_wenable,
  input ram_w16_l512_id19_1_0_enable,
  input [8-1:0] ram_w16_l512_id19_1_1_addr,
  output [16-1:0] ram_w16_l512_id19_1_1_rdata,
  input [16-1:0] ram_w16_l512_id19_1_1_wdata,
  input ram_w16_l512_id19_1_1_wenable,
  input ram_w16_l512_id19_1_1_enable
);

  reg [16-1:0] ram_w16_l512_id19_1_0_rdata_out;
  assign ram_w16_l512_id19_1_0_rdata = ram_w16_l512_id19_1_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id19_1_1_rdata_out;
  assign ram_w16_l512_id19_1_1_rdata = ram_w16_l512_id19_1_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id19_1_0_enable) begin
      if(ram_w16_l512_id19_1_0_wenable) begin
        mem[ram_w16_l512_id19_1_0_addr] <= ram_w16_l512_id19_1_0_wdata;
        ram_w16_l512_id19_1_0_rdata_out <= ram_w16_l512_id19_1_0_wdata;
      end else begin
        ram_w16_l512_id19_1_0_rdata_out <= mem[ram_w16_l512_id19_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id19_1_1_enable) begin
      if(ram_w16_l512_id19_1_1_wenable) begin
        mem[ram_w16_l512_id19_1_1_addr] <= ram_w16_l512_id19_1_1_wdata;
        ram_w16_l512_id19_1_1_rdata_out <= ram_w16_l512_id19_1_1_wdata;
      end else begin
        ram_w16_l512_id19_1_1_rdata_out <= mem[ram_w16_l512_id19_1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id20_0
(
  input CLK,
  input [8-1:0] ram_w16_l512_id20_0_0_addr,
  output [16-1:0] ram_w16_l512_id20_0_0_rdata,
  input [16-1:0] ram_w16_l512_id20_0_0_wdata,
  input ram_w16_l512_id20_0_0_wenable,
  input ram_w16_l512_id20_0_0_enable,
  input [8-1:0] ram_w16_l512_id20_0_1_addr,
  output [16-1:0] ram_w16_l512_id20_0_1_rdata,
  input [16-1:0] ram_w16_l512_id20_0_1_wdata,
  input ram_w16_l512_id20_0_1_wenable,
  input ram_w16_l512_id20_0_1_enable
);

  reg [16-1:0] ram_w16_l512_id20_0_0_rdata_out;
  assign ram_w16_l512_id20_0_0_rdata = ram_w16_l512_id20_0_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id20_0_1_rdata_out;
  assign ram_w16_l512_id20_0_1_rdata = ram_w16_l512_id20_0_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id20_0_0_enable) begin
      if(ram_w16_l512_id20_0_0_wenable) begin
        mem[ram_w16_l512_id20_0_0_addr] <= ram_w16_l512_id20_0_0_wdata;
        ram_w16_l512_id20_0_0_rdata_out <= ram_w16_l512_id20_0_0_wdata;
      end else begin
        ram_w16_l512_id20_0_0_rdata_out <= mem[ram_w16_l512_id20_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id20_0_1_enable) begin
      if(ram_w16_l512_id20_0_1_wenable) begin
        mem[ram_w16_l512_id20_0_1_addr] <= ram_w16_l512_id20_0_1_wdata;
        ram_w16_l512_id20_0_1_rdata_out <= ram_w16_l512_id20_0_1_wdata;
      end else begin
        ram_w16_l512_id20_0_1_rdata_out <= mem[ram_w16_l512_id20_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id20_1
(
  input CLK,
  input [8-1:0] ram_w16_l512_id20_1_0_addr,
  output [16-1:0] ram_w16_l512_id20_1_0_rdata,
  input [16-1:0] ram_w16_l512_id20_1_0_wdata,
  input ram_w16_l512_id20_1_0_wenable,
  input ram_w16_l512_id20_1_0_enable,
  input [8-1:0] ram_w16_l512_id20_1_1_addr,
  output [16-1:0] ram_w16_l512_id20_1_1_rdata,
  input [16-1:0] ram_w16_l512_id20_1_1_wdata,
  input ram_w16_l512_id20_1_1_wenable,
  input ram_w16_l512_id20_1_1_enable
);

  reg [16-1:0] ram_w16_l512_id20_1_0_rdata_out;
  assign ram_w16_l512_id20_1_0_rdata = ram_w16_l512_id20_1_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id20_1_1_rdata_out;
  assign ram_w16_l512_id20_1_1_rdata = ram_w16_l512_id20_1_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id20_1_0_enable) begin
      if(ram_w16_l512_id20_1_0_wenable) begin
        mem[ram_w16_l512_id20_1_0_addr] <= ram_w16_l512_id20_1_0_wdata;
        ram_w16_l512_id20_1_0_rdata_out <= ram_w16_l512_id20_1_0_wdata;
      end else begin
        ram_w16_l512_id20_1_0_rdata_out <= mem[ram_w16_l512_id20_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id20_1_1_enable) begin
      if(ram_w16_l512_id20_1_1_wenable) begin
        mem[ram_w16_l512_id20_1_1_addr] <= ram_w16_l512_id20_1_1_wdata;
        ram_w16_l512_id20_1_1_rdata_out <= ram_w16_l512_id20_1_1_wdata;
      end else begin
        ram_w16_l512_id20_1_1_rdata_out <= mem[ram_w16_l512_id20_1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id21_0
(
  input CLK,
  input [8-1:0] ram_w16_l512_id21_0_0_addr,
  output [16-1:0] ram_w16_l512_id21_0_0_rdata,
  input [16-1:0] ram_w16_l512_id21_0_0_wdata,
  input ram_w16_l512_id21_0_0_wenable,
  input ram_w16_l512_id21_0_0_enable,
  input [8-1:0] ram_w16_l512_id21_0_1_addr,
  output [16-1:0] ram_w16_l512_id21_0_1_rdata,
  input [16-1:0] ram_w16_l512_id21_0_1_wdata,
  input ram_w16_l512_id21_0_1_wenable,
  input ram_w16_l512_id21_0_1_enable
);

  reg [16-1:0] ram_w16_l512_id21_0_0_rdata_out;
  assign ram_w16_l512_id21_0_0_rdata = ram_w16_l512_id21_0_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id21_0_1_rdata_out;
  assign ram_w16_l512_id21_0_1_rdata = ram_w16_l512_id21_0_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id21_0_0_enable) begin
      if(ram_w16_l512_id21_0_0_wenable) begin
        mem[ram_w16_l512_id21_0_0_addr] <= ram_w16_l512_id21_0_0_wdata;
        ram_w16_l512_id21_0_0_rdata_out <= ram_w16_l512_id21_0_0_wdata;
      end else begin
        ram_w16_l512_id21_0_0_rdata_out <= mem[ram_w16_l512_id21_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id21_0_1_enable) begin
      if(ram_w16_l512_id21_0_1_wenable) begin
        mem[ram_w16_l512_id21_0_1_addr] <= ram_w16_l512_id21_0_1_wdata;
        ram_w16_l512_id21_0_1_rdata_out <= ram_w16_l512_id21_0_1_wdata;
      end else begin
        ram_w16_l512_id21_0_1_rdata_out <= mem[ram_w16_l512_id21_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id21_1
(
  input CLK,
  input [8-1:0] ram_w16_l512_id21_1_0_addr,
  output [16-1:0] ram_w16_l512_id21_1_0_rdata,
  input [16-1:0] ram_w16_l512_id21_1_0_wdata,
  input ram_w16_l512_id21_1_0_wenable,
  input ram_w16_l512_id21_1_0_enable,
  input [8-1:0] ram_w16_l512_id21_1_1_addr,
  output [16-1:0] ram_w16_l512_id21_1_1_rdata,
  input [16-1:0] ram_w16_l512_id21_1_1_wdata,
  input ram_w16_l512_id21_1_1_wenable,
  input ram_w16_l512_id21_1_1_enable
);

  reg [16-1:0] ram_w16_l512_id21_1_0_rdata_out;
  assign ram_w16_l512_id21_1_0_rdata = ram_w16_l512_id21_1_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id21_1_1_rdata_out;
  assign ram_w16_l512_id21_1_1_rdata = ram_w16_l512_id21_1_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id21_1_0_enable) begin
      if(ram_w16_l512_id21_1_0_wenable) begin
        mem[ram_w16_l512_id21_1_0_addr] <= ram_w16_l512_id21_1_0_wdata;
        ram_w16_l512_id21_1_0_rdata_out <= ram_w16_l512_id21_1_0_wdata;
      end else begin
        ram_w16_l512_id21_1_0_rdata_out <= mem[ram_w16_l512_id21_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id21_1_1_enable) begin
      if(ram_w16_l512_id21_1_1_wenable) begin
        mem[ram_w16_l512_id21_1_1_addr] <= ram_w16_l512_id21_1_1_wdata;
        ram_w16_l512_id21_1_1_rdata_out <= ram_w16_l512_id21_1_1_wdata;
      end else begin
        ram_w16_l512_id21_1_1_rdata_out <= mem[ram_w16_l512_id21_1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id22_0
(
  input CLK,
  input [8-1:0] ram_w16_l512_id22_0_0_addr,
  output [16-1:0] ram_w16_l512_id22_0_0_rdata,
  input [16-1:0] ram_w16_l512_id22_0_0_wdata,
  input ram_w16_l512_id22_0_0_wenable,
  input ram_w16_l512_id22_0_0_enable,
  input [8-1:0] ram_w16_l512_id22_0_1_addr,
  output [16-1:0] ram_w16_l512_id22_0_1_rdata,
  input [16-1:0] ram_w16_l512_id22_0_1_wdata,
  input ram_w16_l512_id22_0_1_wenable,
  input ram_w16_l512_id22_0_1_enable
);

  reg [16-1:0] ram_w16_l512_id22_0_0_rdata_out;
  assign ram_w16_l512_id22_0_0_rdata = ram_w16_l512_id22_0_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id22_0_1_rdata_out;
  assign ram_w16_l512_id22_0_1_rdata = ram_w16_l512_id22_0_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id22_0_0_enable) begin
      if(ram_w16_l512_id22_0_0_wenable) begin
        mem[ram_w16_l512_id22_0_0_addr] <= ram_w16_l512_id22_0_0_wdata;
        ram_w16_l512_id22_0_0_rdata_out <= ram_w16_l512_id22_0_0_wdata;
      end else begin
        ram_w16_l512_id22_0_0_rdata_out <= mem[ram_w16_l512_id22_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id22_0_1_enable) begin
      if(ram_w16_l512_id22_0_1_wenable) begin
        mem[ram_w16_l512_id22_0_1_addr] <= ram_w16_l512_id22_0_1_wdata;
        ram_w16_l512_id22_0_1_rdata_out <= ram_w16_l512_id22_0_1_wdata;
      end else begin
        ram_w16_l512_id22_0_1_rdata_out <= mem[ram_w16_l512_id22_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id22_1
(
  input CLK,
  input [8-1:0] ram_w16_l512_id22_1_0_addr,
  output [16-1:0] ram_w16_l512_id22_1_0_rdata,
  input [16-1:0] ram_w16_l512_id22_1_0_wdata,
  input ram_w16_l512_id22_1_0_wenable,
  input ram_w16_l512_id22_1_0_enable,
  input [8-1:0] ram_w16_l512_id22_1_1_addr,
  output [16-1:0] ram_w16_l512_id22_1_1_rdata,
  input [16-1:0] ram_w16_l512_id22_1_1_wdata,
  input ram_w16_l512_id22_1_1_wenable,
  input ram_w16_l512_id22_1_1_enable
);

  reg [16-1:0] ram_w16_l512_id22_1_0_rdata_out;
  assign ram_w16_l512_id22_1_0_rdata = ram_w16_l512_id22_1_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id22_1_1_rdata_out;
  assign ram_w16_l512_id22_1_1_rdata = ram_w16_l512_id22_1_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id22_1_0_enable) begin
      if(ram_w16_l512_id22_1_0_wenable) begin
        mem[ram_w16_l512_id22_1_0_addr] <= ram_w16_l512_id22_1_0_wdata;
        ram_w16_l512_id22_1_0_rdata_out <= ram_w16_l512_id22_1_0_wdata;
      end else begin
        ram_w16_l512_id22_1_0_rdata_out <= mem[ram_w16_l512_id22_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id22_1_1_enable) begin
      if(ram_w16_l512_id22_1_1_wenable) begin
        mem[ram_w16_l512_id22_1_1_addr] <= ram_w16_l512_id22_1_1_wdata;
        ram_w16_l512_id22_1_1_rdata_out <= ram_w16_l512_id22_1_1_wdata;
      end else begin
        ram_w16_l512_id22_1_1_rdata_out <= mem[ram_w16_l512_id22_1_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id23_0
(
  input CLK,
  input [8-1:0] ram_w16_l512_id23_0_0_addr,
  output [16-1:0] ram_w16_l512_id23_0_0_rdata,
  input [16-1:0] ram_w16_l512_id23_0_0_wdata,
  input ram_w16_l512_id23_0_0_wenable,
  input ram_w16_l512_id23_0_0_enable,
  input [8-1:0] ram_w16_l512_id23_0_1_addr,
  output [16-1:0] ram_w16_l512_id23_0_1_rdata,
  input [16-1:0] ram_w16_l512_id23_0_1_wdata,
  input ram_w16_l512_id23_0_1_wenable,
  input ram_w16_l512_id23_0_1_enable
);

  reg [16-1:0] ram_w16_l512_id23_0_0_rdata_out;
  assign ram_w16_l512_id23_0_0_rdata = ram_w16_l512_id23_0_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id23_0_1_rdata_out;
  assign ram_w16_l512_id23_0_1_rdata = ram_w16_l512_id23_0_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id23_0_0_enable) begin
      if(ram_w16_l512_id23_0_0_wenable) begin
        mem[ram_w16_l512_id23_0_0_addr] <= ram_w16_l512_id23_0_0_wdata;
        ram_w16_l512_id23_0_0_rdata_out <= ram_w16_l512_id23_0_0_wdata;
      end else begin
        ram_w16_l512_id23_0_0_rdata_out <= mem[ram_w16_l512_id23_0_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id23_0_1_enable) begin
      if(ram_w16_l512_id23_0_1_wenable) begin
        mem[ram_w16_l512_id23_0_1_addr] <= ram_w16_l512_id23_0_1_wdata;
        ram_w16_l512_id23_0_1_rdata_out <= ram_w16_l512_id23_0_1_wdata;
      end else begin
        ram_w16_l512_id23_0_1_rdata_out <= mem[ram_w16_l512_id23_0_1_addr];
      end
    end 
  end


endmodule



module ram_w16_l512_id23_1
(
  input CLK,
  input [8-1:0] ram_w16_l512_id23_1_0_addr,
  output [16-1:0] ram_w16_l512_id23_1_0_rdata,
  input [16-1:0] ram_w16_l512_id23_1_0_wdata,
  input ram_w16_l512_id23_1_0_wenable,
  input ram_w16_l512_id23_1_0_enable,
  input [8-1:0] ram_w16_l512_id23_1_1_addr,
  output [16-1:0] ram_w16_l512_id23_1_1_rdata,
  input [16-1:0] ram_w16_l512_id23_1_1_wdata,
  input ram_w16_l512_id23_1_1_wenable,
  input ram_w16_l512_id23_1_1_enable
);

  reg [16-1:0] ram_w16_l512_id23_1_0_rdata_out;
  assign ram_w16_l512_id23_1_0_rdata = ram_w16_l512_id23_1_0_rdata_out;
  reg [16-1:0] ram_w16_l512_id23_1_1_rdata_out;
  assign ram_w16_l512_id23_1_1_rdata = ram_w16_l512_id23_1_1_rdata_out;
  reg [16-1:0] mem [0:256-1];

  always @(posedge CLK) begin
    if(ram_w16_l512_id23_1_0_enable) begin
      if(ram_w16_l512_id23_1_0_wenable) begin
        mem[ram_w16_l512_id23_1_0_addr] <= ram_w16_l512_id23_1_0_wdata;
        ram_w16_l512_id23_1_0_rdata_out <= ram_w16_l512_id23_1_0_wdata;
      end else begin
        ram_w16_l512_id23_1_0_rdata_out <= mem[ram_w16_l512_id23_1_0_addr];
      end
    end 
  end


  always @(posedge CLK) begin
    if(ram_w16_l512_id23_1_1_enable) begin
      if(ram_w16_l512_id23_1_1_wenable) begin
        mem[ram_w16_l512_id23_1_1_addr] <= ram_w16_l512_id23_1_1_wdata;
        ram_w16_l512_id23_1_1_rdata_out <= ram_w16_l512_id23_1_1_wdata;
      end else begin
        ram_w16_l512_id23_1_1_rdata_out <= mem[ram_w16_l512_id23_1_1_addr];
      end
    end 
  end


endmodule



module madd_9
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_9
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_9
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_10
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_10
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_10
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_11
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_11
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_11
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_12
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_12
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_12
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_13
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_13
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_13
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_14
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_14
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_14
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_15
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_15
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_15
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_16
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_16
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_16
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module madd_17
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);


  madd_core_17
  madd
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c),
    .d(d)
  );


endmodule



module madd_core_17
(
  input CLK,
  input update,
  input [16-1:0] a,
  input [16-1:0] b,
  input [16-1:0] c,
  output [32-1:0] d
);

  reg signed [16-1:0] _a;
  reg signed [16-1:0] _b;
  reg signed [16-1:0] _c;
  wire signed [32-1:0] _mul;
  wire signed [32-1:0] _madd;
  reg signed [32-1:0] _pipe_madd0;
  reg signed [32-1:0] _pipe_madd1;
  assign _mul = _a * _b;
  assign _madd = _mul + _c;
  assign d = _pipe_madd1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _c <= c;
      _pipe_madd0 <= _madd;
      _pipe_madd1 <= _pipe_madd0;
    end 
  end


endmodule



module multiplier_1
(
  input CLK,
  input update,
  input [64-1:0] a,
  input [16-1:0] b,
  output [80-1:0] c
);


  multiplier_core_1
  mult
  (
    .CLK(CLK),
    .update(update),
    .a(a),
    .b(b),
    .c(c)
  );


endmodule



module multiplier_core_1
(
  input CLK,
  input update,
  input [64-1:0] a,
  input [16-1:0] b,
  output [80-1:0] c
);

  reg signed [64-1:0] _a;
  reg signed [16-1:0] _b;
  wire signed [80-1:0] _mul;
  reg signed [80-1:0] _pipe_mul0;
  reg signed [80-1:0] _pipe_mul1;
  assign _mul = _a * _b;
  assign c = _pipe_mul1;

  always @(posedge CLK) begin
    if(update) begin
      _a <= a;
      _b <= b;
      _pipe_mul0 <= _mul;
      _pipe_mul1 <= _pipe_mul0;
    end 
  end


endmodule

